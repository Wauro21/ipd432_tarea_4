`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 01/06/2022 11:35:51 PM
// Design Name:
// Module Name: op_module
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
// Instantation template
/*------------------------------------------
op_module #(
  .N_INPUTS(),
  .I_WIDTH()
)
OP_MOD
(
  .cmd(),
  .enable(),
  .bram_sel(),
  .A(),
  .B(),
  .out()
);
------------------------------------------*/

module op_module#(
  parameter N_INPUTS = 1024,
  parameter I_WIDTH = 8,
  parameter CMD_WIDTH = 3,
  parameter CYCLES_WAIT = 11
  )
  (
  	input logic clk,
  	input logic reset,
    input logic [CMD_WIDTH-1:0] cmd,
    input logic enable,
    input logic bram_sel,
    input logic [N_INPUTS-1:0][I_WIDTH-1:0] A,
    input logic [N_INPUTS-1:0][I_WIDTH-1:0] B,
    output logic [I_WIDTH*3-1:0] out,
	output logic op_done
  );

  eucDis_0 EUC_HLS (
  .C_ap_vld(op_done),  // output wire C_ap_vld
  .ap_clk(clk),      // input wire ap_clk
  .ap_rst(reset),      // input wire ap_rst
  .ap_start(enable),  // input wire ap_start
  .ap_done(),    // output wire ap_done
  .ap_idle(),    // output wire ap_idle
  .ap_ready(),  // output wire ap_ready
  .A_0(A[0]),            // input wire [7 : 0] A_0
  .A_1(A[1]),            // input wire [7 : 0] A_1
  .A_2(A[2]),            // input wire [7 : 0] A_2
  .A_3(A[3]),            // input wire [7 : 0] A_3
  .A_4(A[4]),            // input wire [7 : 0] A_4
  .A_5(A[5]),            // input wire [7 : 0] A_5
  .A_6(A[6]),            // input wire [7 : 0] A_6
  .A_7(A[7]),            // input wire [7 : 0] A_7
  .A_8(A[8]),            // input wire [7 : 0] A_8
  .A_9(A[9]),            // input wire [7 : 0] A_9
  .A_10(A[10]),          // input wire [7 : 0] A_10
  .A_11(A[11]),          // input wire [7 : 0] A_11
  .A_12(A[12]),          // input wire [7 : 0] A_12
  .A_13(A[13]),          // input wire [7 : 0] A_13
  .A_14(A[14]),          // input wire [7 : 0] A_14
  .A_15(A[15]),          // input wire [7 : 0] A_15
  .A_16(A[16]),          // input wire [7 : 0] A_16
  .A_17(A[17]),          // input wire [7 : 0] A_17
  .A_18(A[18]),          // input wire [7 : 0] A_18
  .A_19(A[19]),          // input wire [7 : 0] A_19
  .A_20(A[20]),          // input wire [7 : 0] A_20
  .A_21(A[21]),          // input wire [7 : 0] A_21
  .A_22(A[22]),          // input wire [7 : 0] A_22
  .A_23(A[23]),          // input wire [7 : 0] A_23
  .A_24(A[24]),          // input wire [7 : 0] A_24
  .A_25(A[25]),          // input wire [7 : 0] A_25
  .A_26(A[26]),          // input wire [7 : 0] A_26
  .A_27(A[27]),          // input wire [7 : 0] A_27
  .A_28(A[28]),          // input wire [7 : 0] A_28
  .A_29(A[29]),          // input wire [7 : 0] A_29
  .A_30(A[30]),          // input wire [7 : 0] A_30
  .A_31(A[31]),          // input wire [7 : 0] A_31
  .A_32(A[32]),          // input wire [7 : 0] A_32
  .A_33(A[33]),          // input wire [7 : 0] A_33
  .A_34(A[34]),          // input wire [7 : 0] A_34
  .A_35(A[35]),          // input wire [7 : 0] A_35
  .A_36(A[36]),          // input wire [7 : 0] A_36
  .A_37(A[37]),          // input wire [7 : 0] A_37
  .A_38(A[38]),          // input wire [7 : 0] A_38
  .A_39(A[39]),          // input wire [7 : 0] A_39
  .A_40(A[40]),          // input wire [7 : 0] A_40
  .A_41(A[41]),          // input wire [7 : 0] A_41
  .A_42(A[42]),          // input wire [7 : 0] A_42
  .A_43(A[43]),          // input wire [7 : 0] A_43
  .A_44(A[44]),          // input wire [7 : 0] A_44
  .A_45(A[45]),          // input wire [7 : 0] A_45
  .A_46(A[46]),          // input wire [7 : 0] A_46
  .A_47(A[47]),          // input wire [7 : 0] A_47
  .A_48(A[48]),          // input wire [7 : 0] A_48
  .A_49(A[49]),          // input wire [7 : 0] A_49
  .A_50(A[50]),          // input wire [7 : 0] A_50
  .A_51(A[51]),          // input wire [7 : 0] A_51
  .A_52(A[52]),          // input wire [7 : 0] A_52
  .A_53(A[53]),          // input wire [7 : 0] A_53
  .A_54(A[54]),          // input wire [7 : 0] A_54
  .A_55(A[55]),          // input wire [7 : 0] A_55
  .A_56(A[56]),          // input wire [7 : 0] A_56
  .A_57(A[57]),          // input wire [7 : 0] A_57
  .A_58(A[58]),          // input wire [7 : 0] A_58
  .A_59(A[59]),          // input wire [7 : 0] A_59
  .A_60(A[60]),          // input wire [7 : 0] A_60
  .A_61(A[61]),          // input wire [7 : 0] A_61
  .A_62(A[62]),          // input wire [7 : 0] A_62
  .A_63(A[63]),          // input wire [7 : 0] A_63
  .A_64(A[64]),          // input wire [7 : 0] A_64
  .A_65(A[65]),          // input wire [7 : 0] A_65
  .A_66(A[66]),          // input wire [7 : 0] A_66
  .A_67(A[67]),          // input wire [7 : 0] A_67
  .A_68(A[68]),          // input wire [7 : 0] A_68
  .A_69(A[69]),          // input wire [7 : 0] A_69
  .A_70(A[70]),          // input wire [7 : 0] A_70
  .A_71(A[71]),          // input wire [7 : 0] A_71
  .A_72(A[72]),          // input wire [7 : 0] A_72
  .A_73(A[73]),          // input wire [7 : 0] A_73
  .A_74(A[74]),          // input wire [7 : 0] A_74
  .A_75(A[75]),          // input wire [7 : 0] A_75
  .A_76(A[76]),          // input wire [7 : 0] A_76
  .A_77(A[77]),          // input wire [7 : 0] A_77
  .A_78(A[78]),          // input wire [7 : 0] A_78
  .A_79(A[79]),          // input wire [7 : 0] A_79
  .A_80(A[80]),          // input wire [7 : 0] A_80
  .A_81(A[81]),          // input wire [7 : 0] A_81
  .A_82(A[82]),          // input wire [7 : 0] A_82
  .A_83(A[83]),          // input wire [7 : 0] A_83
  .A_84(A[84]),          // input wire [7 : 0] A_84
  .A_85(A[85]),          // input wire [7 : 0] A_85
  .A_86(A[86]),          // input wire [7 : 0] A_86
  .A_87(A[87]),          // input wire [7 : 0] A_87
  .A_88(A[88]),          // input wire [7 : 0] A_88
  .A_89(A[89]),          // input wire [7 : 0] A_89
  .A_90(A[90]),          // input wire [7 : 0] A_90
  .A_91(A[91]),          // input wire [7 : 0] A_91
  .A_92(A[92]),          // input wire [7 : 0] A_92
  .A_93(A[93]),          // input wire [7 : 0] A_93
  .A_94(A[94]),          // input wire [7 : 0] A_94
  .A_95(A[95]),          // input wire [7 : 0] A_95
  .A_96(A[96]),          // input wire [7 : 0] A_96
  .A_97(A[97]),          // input wire [7 : 0] A_97
  .A_98(A[98]),          // input wire [7 : 0] A_98
  .A_99(A[99]),          // input wire [7 : 0] A_99
  .A_100(A[100]),        // input wire [7 : 0] A_100
  .A_101(A[101]),        // input wire [7 : 0] A_101
  .A_102(A[102]),        // input wire [7 : 0] A_102
  .A_103(A[103]),        // input wire [7 : 0] A_103
  .A_104(A[104]),        // input wire [7 : 0] A_104
  .A_105(A[105]),        // input wire [7 : 0] A_105
  .A_106(A[106]),        // input wire [7 : 0] A_106
  .A_107(A[107]),        // input wire [7 : 0] A_107
  .A_108(A[108]),        // input wire [7 : 0] A_108
  .A_109(A[109]),        // input wire [7 : 0] A_109
  .A_110(A[110]),        // input wire [7 : 0] A_110
  .A_111(A[111]),        // input wire [7 : 0] A_111
  .A_112(A[112]),        // input wire [7 : 0] A_112
  .A_113(A[113]),        // input wire [7 : 0] A_113
  .A_114(A[114]),        // input wire [7 : 0] A_114
  .A_115(A[115]),        // input wire [7 : 0] A_115
  .A_116(A[116]),        // input wire [7 : 0] A_116
  .A_117(A[117]),        // input wire [7 : 0] A_117
  .A_118(A[118]),        // input wire [7 : 0] A_118
  .A_119(A[119]),        // input wire [7 : 0] A_119
  .A_120(A[120]),        // input wire [7 : 0] A_120
  .A_121(A[121]),        // input wire [7 : 0] A_121
  .A_122(A[122]),        // input wire [7 : 0] A_122
  .A_123(A[123]),        // input wire [7 : 0] A_123
  .A_124(A[124]),        // input wire [7 : 0] A_124
  .A_125(A[125]),        // input wire [7 : 0] A_125
  .A_126(A[126]),        // input wire [7 : 0] A_126
  .A_127(A[127]),        // input wire [7 : 0] A_127
  .A_128(A[128]),        // input wire [7 : 0] A_128
  .A_129(A[129]),        // input wire [7 : 0] A_129
  .A_130(A[130]),        // input wire [7 : 0] A_130
  .A_131(A[131]),        // input wire [7 : 0] A_131
  .A_132(A[132]),        // input wire [7 : 0] A_132
  .A_133(A[133]),        // input wire [7 : 0] A_133
  .A_134(A[134]),        // input wire [7 : 0] A_134
  .A_135(A[135]),        // input wire [7 : 0] A_135
  .A_136(A[136]),        // input wire [7 : 0] A_136
  .A_137(A[137]),        // input wire [7 : 0] A_137
  .A_138(A[138]),        // input wire [7 : 0] A_138
  .A_139(A[139]),        // input wire [7 : 0] A_139
  .A_140(A[140]),        // input wire [7 : 0] A_140
  .A_141(A[141]),        // input wire [7 : 0] A_141
  .A_142(A[142]),        // input wire [7 : 0] A_142
  .A_143(A[143]),        // input wire [7 : 0] A_143
  .A_144(A[144]),        // input wire [7 : 0] A_144
  .A_145(A[145]),        // input wire [7 : 0] A_145
  .A_146(A[146]),        // input wire [7 : 0] A_146
  .A_147(A[147]),        // input wire [7 : 0] A_147
  .A_148(A[148]),        // input wire [7 : 0] A_148
  .A_149(A[149]),        // input wire [7 : 0] A_149
  .A_150(A[150]),        // input wire [7 : 0] A_150
  .A_151(A[151]),        // input wire [7 : 0] A_151
  .A_152(A[152]),        // input wire [7 : 0] A_152
  .A_153(A[153]),        // input wire [7 : 0] A_153
  .A_154(A[154]),        // input wire [7 : 0] A_154
  .A_155(A[155]),        // input wire [7 : 0] A_155
  .A_156(A[156]),        // input wire [7 : 0] A_156
  .A_157(A[157]),        // input wire [7 : 0] A_157
  .A_158(A[158]),        // input wire [7 : 0] A_158
  .A_159(A[159]),        // input wire [7 : 0] A_159
  .A_160(A[160]),        // input wire [7 : 0] A_160
  .A_161(A[161]),        // input wire [7 : 0] A_161
  .A_162(A[162]),        // input wire [7 : 0] A_162
  .A_163(A[163]),        // input wire [7 : 0] A_163
  .A_164(A[164]),        // input wire [7 : 0] A_164
  .A_165(A[165]),        // input wire [7 : 0] A_165
  .A_166(A[166]),        // input wire [7 : 0] A_166
  .A_167(A[167]),        // input wire [7 : 0] A_167
  .A_168(A[168]),        // input wire [7 : 0] A_168
  .A_169(A[169]),        // input wire [7 : 0] A_169
  .A_170(A[170]),        // input wire [7 : 0] A_170
  .A_171(A[171]),        // input wire [7 : 0] A_171
  .A_172(A[172]),        // input wire [7 : 0] A_172
  .A_173(A[173]),        // input wire [7 : 0] A_173
  .A_174(A[174]),        // input wire [7 : 0] A_174
  .A_175(A[175]),        // input wire [7 : 0] A_175
  .A_176(A[176]),        // input wire [7 : 0] A_176
  .A_177(A[177]),        // input wire [7 : 0] A_177
  .A_178(A[178]),        // input wire [7 : 0] A_178
  .A_179(A[179]),        // input wire [7 : 0] A_179
  .A_180(A[180]),        // input wire [7 : 0] A_180
  .A_181(A[181]),        // input wire [7 : 0] A_181
  .A_182(A[182]),        // input wire [7 : 0] A_182
  .A_183(A[183]),        // input wire [7 : 0] A_183
  .A_184(A[184]),        // input wire [7 : 0] A_184
  .A_185(A[185]),        // input wire [7 : 0] A_185
  .A_186(A[186]),        // input wire [7 : 0] A_186
  .A_187(A[187]),        // input wire [7 : 0] A_187
  .A_188(A[188]),        // input wire [7 : 0] A_188
  .A_189(A[189]),        // input wire [7 : 0] A_189
  .A_190(A[190]),        // input wire [7 : 0] A_190
  .A_191(A[191]),        // input wire [7 : 0] A_191
  .A_192(A[192]),        // input wire [7 : 0] A_192
  .A_193(A[193]),        // input wire [7 : 0] A_193
  .A_194(A[194]),        // input wire [7 : 0] A_194
  .A_195(A[195]),        // input wire [7 : 0] A_195
  .A_196(A[196]),        // input wire [7 : 0] A_196
  .A_197(A[197]),        // input wire [7 : 0] A_197
  .A_198(A[198]),        // input wire [7 : 0] A_198
  .A_199(A[199]),        // input wire [7 : 0] A_199
  .A_200(A[200]),        // input wire [7 : 0] A_200
  .A_201(A[201]),        // input wire [7 : 0] A_201
  .A_202(A[202]),        // input wire [7 : 0] A_202
  .A_203(A[203]),        // input wire [7 : 0] A_203
  .A_204(A[204]),        // input wire [7 : 0] A_204
  .A_205(A[205]),        // input wire [7 : 0] A_205
  .A_206(A[206]),        // input wire [7 : 0] A_206
  .A_207(A[207]),        // input wire [7 : 0] A_207
  .A_208(A[208]),        // input wire [7 : 0] A_208
  .A_209(A[209]),        // input wire [7 : 0] A_209
  .A_210(A[210]),        // input wire [7 : 0] A_210
  .A_211(A[211]),        // input wire [7 : 0] A_211
  .A_212(A[212]),        // input wire [7 : 0] A_212
  .A_213(A[213]),        // input wire [7 : 0] A_213
  .A_214(A[214]),        // input wire [7 : 0] A_214
  .A_215(A[215]),        // input wire [7 : 0] A_215
  .A_216(A[216]),        // input wire [7 : 0] A_216
  .A_217(A[217]),        // input wire [7 : 0] A_217
  .A_218(A[218]),        // input wire [7 : 0] A_218
  .A_219(A[219]),        // input wire [7 : 0] A_219
  .A_220(A[220]),        // input wire [7 : 0] A_220
  .A_221(A[221]),        // input wire [7 : 0] A_221
  .A_222(A[222]),        // input wire [7 : 0] A_222
  .A_223(A[223]),        // input wire [7 : 0] A_223
  .A_224(A[224]),        // input wire [7 : 0] A_224
  .A_225(A[225]),        // input wire [7 : 0] A_225
  .A_226(A[226]),        // input wire [7 : 0] A_226
  .A_227(A[227]),        // input wire [7 : 0] A_227
  .A_228(A[228]),        // input wire [7 : 0] A_228
  .A_229(A[229]),        // input wire [7 : 0] A_229
  .A_230(A[230]),        // input wire [7 : 0] A_230
  .A_231(A[231]),        // input wire [7 : 0] A_231
  .A_232(A[232]),        // input wire [7 : 0] A_232
  .A_233(A[233]),        // input wire [7 : 0] A_233
  .A_234(A[234]),        // input wire [7 : 0] A_234
  .A_235(A[235]),        // input wire [7 : 0] A_235
  .A_236(A[236]),        // input wire [7 : 0] A_236
  .A_237(A[237]),        // input wire [7 : 0] A_237
  .A_238(A[238]),        // input wire [7 : 0] A_238
  .A_239(A[239]),        // input wire [7 : 0] A_239
  .A_240(A[240]),        // input wire [7 : 0] A_240
  .A_241(A[241]),        // input wire [7 : 0] A_241
  .A_242(A[242]),        // input wire [7 : 0] A_242
  .A_243(A[243]),        // input wire [7 : 0] A_243
  .A_244(A[244]),        // input wire [7 : 0] A_244
  .A_245(A[245]),        // input wire [7 : 0] A_245
  .A_246(A[246]),        // input wire [7 : 0] A_246
  .A_247(A[247]),        // input wire [7 : 0] A_247
  .A_248(A[248]),        // input wire [7 : 0] A_248
  .A_249(A[249]),        // input wire [7 : 0] A_249
  .A_250(A[250]),        // input wire [7 : 0] A_250
  .A_251(A[251]),        // input wire [7 : 0] A_251
  .A_252(A[252]),        // input wire [7 : 0] A_252
  .A_253(A[253]),        // input wire [7 : 0] A_253
  .A_254(A[254]),        // input wire [7 : 0] A_254
  .A_255(A[255]),        // input wire [7 : 0] A_255
  .A_256(A[256]),        // input wire [7 : 0] A_256
  .A_257(A[257]),        // input wire [7 : 0] A_257
  .A_258(A[258]),        // input wire [7 : 0] A_258
  .A_259(A[259]),        // input wire [7 : 0] A_259
  .A_260(A[260]),        // input wire [7 : 0] A_260
  .A_261(A[261]),        // input wire [7 : 0] A_261
  .A_262(A[262]),        // input wire [7 : 0] A_262
  .A_263(A[263]),        // input wire [7 : 0] A_263
  .A_264(A[264]),        // input wire [7 : 0] A_264
  .A_265(A[265]),        // input wire [7 : 0] A_265
  .A_266(A[266]),        // input wire [7 : 0] A_266
  .A_267(A[267]),        // input wire [7 : 0] A_267
  .A_268(A[268]),        // input wire [7 : 0] A_268
  .A_269(A[269]),        // input wire [7 : 0] A_269
  .A_270(A[270]),        // input wire [7 : 0] A_270
  .A_271(A[271]),        // input wire [7 : 0] A_271
  .A_272(A[272]),        // input wire [7 : 0] A_272
  .A_273(A[273]),        // input wire [7 : 0] A_273
  .A_274(A[274]),        // input wire [7 : 0] A_274
  .A_275(A[275]),        // input wire [7 : 0] A_275
  .A_276(A[276]),        // input wire [7 : 0] A_276
  .A_277(A[277]),        // input wire [7 : 0] A_277
  .A_278(A[278]),        // input wire [7 : 0] A_278
  .A_279(A[279]),        // input wire [7 : 0] A_279
  .A_280(A[280]),        // input wire [7 : 0] A_280
  .A_281(A[281]),        // input wire [7 : 0] A_281
  .A_282(A[282]),        // input wire [7 : 0] A_282
  .A_283(A[283]),        // input wire [7 : 0] A_283
  .A_284(A[284]),        // input wire [7 : 0] A_284
  .A_285(A[285]),        // input wire [7 : 0] A_285
  .A_286(A[286]),        // input wire [7 : 0] A_286
  .A_287(A[287]),        // input wire [7 : 0] A_287
  .A_288(A[288]),        // input wire [7 : 0] A_288
  .A_289(A[289]),        // input wire [7 : 0] A_289
  .A_290(A[290]),        // input wire [7 : 0] A_290
  .A_291(A[291]),        // input wire [7 : 0] A_291
  .A_292(A[292]),        // input wire [7 : 0] A_292
  .A_293(A[293]),        // input wire [7 : 0] A_293
  .A_294(A[294]),        // input wire [7 : 0] A_294
  .A_295(A[295]),        // input wire [7 : 0] A_295
  .A_296(A[296]),        // input wire [7 : 0] A_296
  .A_297(A[297]),        // input wire [7 : 0] A_297
  .A_298(A[298]),        // input wire [7 : 0] A_298
  .A_299(A[299]),        // input wire [7 : 0] A_299
  .A_300(A[300]),        // input wire [7 : 0] A_300
  .A_301(A[301]),        // input wire [7 : 0] A_301
  .A_302(A[302]),        // input wire [7 : 0] A_302
  .A_303(A[303]),        // input wire [7 : 0] A_303
  .A_304(A[304]),        // input wire [7 : 0] A_304
  .A_305(A[305]),        // input wire [7 : 0] A_305
  .A_306(A[306]),        // input wire [7 : 0] A_306
  .A_307(A[307]),        // input wire [7 : 0] A_307
  .A_308(A[308]),        // input wire [7 : 0] A_308
  .A_309(A[309]),        // input wire [7 : 0] A_309
  .A_310(A[310]),        // input wire [7 : 0] A_310
  .A_311(A[311]),        // input wire [7 : 0] A_311
  .A_312(A[312]),        // input wire [7 : 0] A_312
  .A_313(A[313]),        // input wire [7 : 0] A_313
  .A_314(A[314]),        // input wire [7 : 0] A_314
  .A_315(A[315]),        // input wire [7 : 0] A_315
  .A_316(A[316]),        // input wire [7 : 0] A_316
  .A_317(A[317]),        // input wire [7 : 0] A_317
  .A_318(A[318]),        // input wire [7 : 0] A_318
  .A_319(A[319]),        // input wire [7 : 0] A_319
  .A_320(A[320]),        // input wire [7 : 0] A_320
  .A_321(A[321]),        // input wire [7 : 0] A_321
  .A_322(A[322]),        // input wire [7 : 0] A_322
  .A_323(A[323]),        // input wire [7 : 0] A_323
  .A_324(A[324]),        // input wire [7 : 0] A_324
  .A_325(A[325]),        // input wire [7 : 0] A_325
  .A_326(A[326]),        // input wire [7 : 0] A_326
  .A_327(A[327]),        // input wire [7 : 0] A_327
  .A_328(A[328]),        // input wire [7 : 0] A_328
  .A_329(A[329]),        // input wire [7 : 0] A_329
  .A_330(A[330]),        // input wire [7 : 0] A_330
  .A_331(A[331]),        // input wire [7 : 0] A_331
  .A_332(A[332]),        // input wire [7 : 0] A_332
  .A_333(A[333]),        // input wire [7 : 0] A_333
  .A_334(A[334]),        // input wire [7 : 0] A_334
  .A_335(A[335]),        // input wire [7 : 0] A_335
  .A_336(A[336]),        // input wire [7 : 0] A_336
  .A_337(A[337]),        // input wire [7 : 0] A_337
  .A_338(A[338]),        // input wire [7 : 0] A_338
  .A_339(A[339]),        // input wire [7 : 0] A_339
  .A_340(A[340]),        // input wire [7 : 0] A_340
  .A_341(A[341]),        // input wire [7 : 0] A_341
  .A_342(A[342]),        // input wire [7 : 0] A_342
  .A_343(A[343]),        // input wire [7 : 0] A_343
  .A_344(A[344]),        // input wire [7 : 0] A_344
  .A_345(A[345]),        // input wire [7 : 0] A_345
  .A_346(A[346]),        // input wire [7 : 0] A_346
  .A_347(A[347]),        // input wire [7 : 0] A_347
  .A_348(A[348]),        // input wire [7 : 0] A_348
  .A_349(A[349]),        // input wire [7 : 0] A_349
  .A_350(A[350]),        // input wire [7 : 0] A_350
  .A_351(A[351]),        // input wire [7 : 0] A_351
  .A_352(A[352]),        // input wire [7 : 0] A_352
  .A_353(A[353]),        // input wire [7 : 0] A_353
  .A_354(A[354]),        // input wire [7 : 0] A_354
  .A_355(A[355]),        // input wire [7 : 0] A_355
  .A_356(A[356]),        // input wire [7 : 0] A_356
  .A_357(A[357]),        // input wire [7 : 0] A_357
  .A_358(A[358]),        // input wire [7 : 0] A_358
  .A_359(A[359]),        // input wire [7 : 0] A_359
  .A_360(A[360]),        // input wire [7 : 0] A_360
  .A_361(A[361]),        // input wire [7 : 0] A_361
  .A_362(A[362]),        // input wire [7 : 0] A_362
  .A_363(A[363]),        // input wire [7 : 0] A_363
  .A_364(A[364]),        // input wire [7 : 0] A_364
  .A_365(A[365]),        // input wire [7 : 0] A_365
  .A_366(A[366]),        // input wire [7 : 0] A_366
  .A_367(A[367]),        // input wire [7 : 0] A_367
  .A_368(A[368]),        // input wire [7 : 0] A_368
  .A_369(A[369]),        // input wire [7 : 0] A_369
  .A_370(A[370]),        // input wire [7 : 0] A_370
  .A_371(A[371]),        // input wire [7 : 0] A_371
  .A_372(A[372]),        // input wire [7 : 0] A_372
  .A_373(A[373]),        // input wire [7 : 0] A_373
  .A_374(A[374]),        // input wire [7 : 0] A_374
  .A_375(A[375]),        // input wire [7 : 0] A_375
  .A_376(A[376]),        // input wire [7 : 0] A_376
  .A_377(A[377]),        // input wire [7 : 0] A_377
  .A_378(A[378]),        // input wire [7 : 0] A_378
  .A_379(A[379]),        // input wire [7 : 0] A_379
  .A_380(A[380]),        // input wire [7 : 0] A_380
  .A_381(A[381]),        // input wire [7 : 0] A_381
  .A_382(A[382]),        // input wire [7 : 0] A_382
  .A_383(A[383]),        // input wire [7 : 0] A_383
  .A_384(A[384]),        // input wire [7 : 0] A_384
  .A_385(A[385]),        // input wire [7 : 0] A_385
  .A_386(A[386]),        // input wire [7 : 0] A_386
  .A_387(A[387]),        // input wire [7 : 0] A_387
  .A_388(A[388]),        // input wire [7 : 0] A_388
  .A_389(A[389]),        // input wire [7 : 0] A_389
  .A_390(A[390]),        // input wire [7 : 0] A_390
  .A_391(A[391]),        // input wire [7 : 0] A_391
  .A_392(A[392]),        // input wire [7 : 0] A_392
  .A_393(A[393]),        // input wire [7 : 0] A_393
  .A_394(A[394]),        // input wire [7 : 0] A_394
  .A_395(A[395]),        // input wire [7 : 0] A_395
  .A_396(A[396]),        // input wire [7 : 0] A_396
  .A_397(A[397]),        // input wire [7 : 0] A_397
  .A_398(A[398]),        // input wire [7 : 0] A_398
  .A_399(A[399]),        // input wire [7 : 0] A_399
  .A_400(A[400]),        // input wire [7 : 0] A_400
  .A_401(A[401]),        // input wire [7 : 0] A_401
  .A_402(A[402]),        // input wire [7 : 0] A_402
  .A_403(A[403]),        // input wire [7 : 0] A_403
  .A_404(A[404]),        // input wire [7 : 0] A_404
  .A_405(A[405]),        // input wire [7 : 0] A_405
  .A_406(A[406]),        // input wire [7 : 0] A_406
  .A_407(A[407]),        // input wire [7 : 0] A_407
  .A_408(A[408]),        // input wire [7 : 0] A_408
  .A_409(A[409]),        // input wire [7 : 0] A_409
  .A_410(A[410]),        // input wire [7 : 0] A_410
  .A_411(A[411]),        // input wire [7 : 0] A_411
  .A_412(A[412]),        // input wire [7 : 0] A_412
  .A_413(A[413]),        // input wire [7 : 0] A_413
  .A_414(A[414]),        // input wire [7 : 0] A_414
  .A_415(A[415]),        // input wire [7 : 0] A_415
  .A_416(A[416]),        // input wire [7 : 0] A_416
  .A_417(A[417]),        // input wire [7 : 0] A_417
  .A_418(A[418]),        // input wire [7 : 0] A_418
  .A_419(A[419]),        // input wire [7 : 0] A_419
  .A_420(A[420]),        // input wire [7 : 0] A_420
  .A_421(A[421]),        // input wire [7 : 0] A_421
  .A_422(A[422]),        // input wire [7 : 0] A_422
  .A_423(A[423]),        // input wire [7 : 0] A_423
  .A_424(A[424]),        // input wire [7 : 0] A_424
  .A_425(A[425]),        // input wire [7 : 0] A_425
  .A_426(A[426]),        // input wire [7 : 0] A_426
  .A_427(A[427]),        // input wire [7 : 0] A_427
  .A_428(A[428]),        // input wire [7 : 0] A_428
  .A_429(A[429]),        // input wire [7 : 0] A_429
  .A_430(A[430]),        // input wire [7 : 0] A_430
  .A_431(A[431]),        // input wire [7 : 0] A_431
  .A_432(A[432]),        // input wire [7 : 0] A_432
  .A_433(A[433]),        // input wire [7 : 0] A_433
  .A_434(A[434]),        // input wire [7 : 0] A_434
  .A_435(A[435]),        // input wire [7 : 0] A_435
  .A_436(A[436]),        // input wire [7 : 0] A_436
  .A_437(A[437]),        // input wire [7 : 0] A_437
  .A_438(A[438]),        // input wire [7 : 0] A_438
  .A_439(A[439]),        // input wire [7 : 0] A_439
  .A_440(A[440]),        // input wire [7 : 0] A_440
  .A_441(A[441]),        // input wire [7 : 0] A_441
  .A_442(A[442]),        // input wire [7 : 0] A_442
  .A_443(A[443]),        // input wire [7 : 0] A_443
  .A_444(A[444]),        // input wire [7 : 0] A_444
  .A_445(A[445]),        // input wire [7 : 0] A_445
  .A_446(A[446]),        // input wire [7 : 0] A_446
  .A_447(A[447]),        // input wire [7 : 0] A_447
  .A_448(A[448]),        // input wire [7 : 0] A_448
  .A_449(A[449]),        // input wire [7 : 0] A_449
  .A_450(A[450]),        // input wire [7 : 0] A_450
  .A_451(A[451]),        // input wire [7 : 0] A_451
  .A_452(A[452]),        // input wire [7 : 0] A_452
  .A_453(A[453]),        // input wire [7 : 0] A_453
  .A_454(A[454]),        // input wire [7 : 0] A_454
  .A_455(A[455]),        // input wire [7 : 0] A_455
  .A_456(A[456]),        // input wire [7 : 0] A_456
  .A_457(A[457]),        // input wire [7 : 0] A_457
  .A_458(A[458]),        // input wire [7 : 0] A_458
  .A_459(A[459]),        // input wire [7 : 0] A_459
  .A_460(A[460]),        // input wire [7 : 0] A_460
  .A_461(A[461]),        // input wire [7 : 0] A_461
  .A_462(A[462]),        // input wire [7 : 0] A_462
  .A_463(A[463]),        // input wire [7 : 0] A_463
  .A_464(A[464]),        // input wire [7 : 0] A_464
  .A_465(A[465]),        // input wire [7 : 0] A_465
  .A_466(A[466]),        // input wire [7 : 0] A_466
  .A_467(A[467]),        // input wire [7 : 0] A_467
  .A_468(A[468]),        // input wire [7 : 0] A_468
  .A_469(A[469]),        // input wire [7 : 0] A_469
  .A_470(A[470]),        // input wire [7 : 0] A_470
  .A_471(A[471]),        // input wire [7 : 0] A_471
  .A_472(A[472]),        // input wire [7 : 0] A_472
  .A_473(A[473]),        // input wire [7 : 0] A_473
  .A_474(A[474]),        // input wire [7 : 0] A_474
  .A_475(A[475]),        // input wire [7 : 0] A_475
  .A_476(A[476]),        // input wire [7 : 0] A_476
  .A_477(A[477]),        // input wire [7 : 0] A_477
  .A_478(A[478]),        // input wire [7 : 0] A_478
  .A_479(A[479]),        // input wire [7 : 0] A_479
  .A_480(A[480]),        // input wire [7 : 0] A_480
  .A_481(A[481]),        // input wire [7 : 0] A_481
  .A_482(A[482]),        // input wire [7 : 0] A_482
  .A_483(A[483]),        // input wire [7 : 0] A_483
  .A_484(A[484]),        // input wire [7 : 0] A_484
  .A_485(A[485]),        // input wire [7 : 0] A_485
  .A_486(A[486]),        // input wire [7 : 0] A_486
  .A_487(A[487]),        // input wire [7 : 0] A_487
  .A_488(A[488]),        // input wire [7 : 0] A_488
  .A_489(A[489]),        // input wire [7 : 0] A_489
  .A_490(A[490]),        // input wire [7 : 0] A_490
  .A_491(A[491]),        // input wire [7 : 0] A_491
  .A_492(A[492]),        // input wire [7 : 0] A_492
  .A_493(A[493]),        // input wire [7 : 0] A_493
  .A_494(A[494]),        // input wire [7 : 0] A_494
  .A_495(A[495]),        // input wire [7 : 0] A_495
  .A_496(A[496]),        // input wire [7 : 0] A_496
  .A_497(A[497]),        // input wire [7 : 0] A_497
  .A_498(A[498]),        // input wire [7 : 0] A_498
  .A_499(A[499]),        // input wire [7 : 0] A_499
  .A_500(A[500]),        // input wire [7 : 0] A_500
  .A_501(A[501]),        // input wire [7 : 0] A_501
  .A_502(A[502]),        // input wire [7 : 0] A_502
  .A_503(A[503]),        // input wire [7 : 0] A_503
  .A_504(A[504]),        // input wire [7 : 0] A_504
  .A_505(A[505]),        // input wire [7 : 0] A_505
  .A_506(A[506]),        // input wire [7 : 0] A_506
  .A_507(A[507]),        // input wire [7 : 0] A_507
  .A_508(A[508]),        // input wire [7 : 0] A_508
  .A_509(A[509]),        // input wire [7 : 0] A_509
  .A_510(A[510]),        // input wire [7 : 0] A_510
  .A_511(A[511]),        // input wire [7 : 0] A_511
  .A_512(A[512]),        // input wire [7 : 0] A_512
  .A_513(A[513]),        // input wire [7 : 0] A_513
  .A_514(A[514]),        // input wire [7 : 0] A_514
  .A_515(A[515]),        // input wire [7 : 0] A_515
  .A_516(A[516]),        // input wire [7 : 0] A_516
  .A_517(A[517]),        // input wire [7 : 0] A_517
  .A_518(A[518]),        // input wire [7 : 0] A_518
  .A_519(A[519]),        // input wire [7 : 0] A_519
  .A_520(A[520]),        // input wire [7 : 0] A_520
  .A_521(A[521]),        // input wire [7 : 0] A_521
  .A_522(A[522]),        // input wire [7 : 0] A_522
  .A_523(A[523]),        // input wire [7 : 0] A_523
  .A_524(A[524]),        // input wire [7 : 0] A_524
  .A_525(A[525]),        // input wire [7 : 0] A_525
  .A_526(A[526]),        // input wire [7 : 0] A_526
  .A_527(A[527]),        // input wire [7 : 0] A_527
  .A_528(A[528]),        // input wire [7 : 0] A_528
  .A_529(A[529]),        // input wire [7 : 0] A_529
  .A_530(A[530]),        // input wire [7 : 0] A_530
  .A_531(A[531]),        // input wire [7 : 0] A_531
  .A_532(A[532]),        // input wire [7 : 0] A_532
  .A_533(A[533]),        // input wire [7 : 0] A_533
  .A_534(A[534]),        // input wire [7 : 0] A_534
  .A_535(A[535]),        // input wire [7 : 0] A_535
  .A_536(A[536]),        // input wire [7 : 0] A_536
  .A_537(A[537]),        // input wire [7 : 0] A_537
  .A_538(A[538]),        // input wire [7 : 0] A_538
  .A_539(A[539]),        // input wire [7 : 0] A_539
  .A_540(A[540]),        // input wire [7 : 0] A_540
  .A_541(A[541]),        // input wire [7 : 0] A_541
  .A_542(A[542]),        // input wire [7 : 0] A_542
  .A_543(A[543]),        // input wire [7 : 0] A_543
  .A_544(A[544]),        // input wire [7 : 0] A_544
  .A_545(A[545]),        // input wire [7 : 0] A_545
  .A_546(A[546]),        // input wire [7 : 0] A_546
  .A_547(A[547]),        // input wire [7 : 0] A_547
  .A_548(A[548]),        // input wire [7 : 0] A_548
  .A_549(A[549]),        // input wire [7 : 0] A_549
  .A_550(A[550]),        // input wire [7 : 0] A_550
  .A_551(A[551]),        // input wire [7 : 0] A_551
  .A_552(A[552]),        // input wire [7 : 0] A_552
  .A_553(A[553]),        // input wire [7 : 0] A_553
  .A_554(A[554]),        // input wire [7 : 0] A_554
  .A_555(A[555]),        // input wire [7 : 0] A_555
  .A_556(A[556]),        // input wire [7 : 0] A_556
  .A_557(A[557]),        // input wire [7 : 0] A_557
  .A_558(A[558]),        // input wire [7 : 0] A_558
  .A_559(A[559]),        // input wire [7 : 0] A_559
  .A_560(A[560]),        // input wire [7 : 0] A_560
  .A_561(A[561]),        // input wire [7 : 0] A_561
  .A_562(A[562]),        // input wire [7 : 0] A_562
  .A_563(A[563]),        // input wire [7 : 0] A_563
  .A_564(A[564]),        // input wire [7 : 0] A_564
  .A_565(A[565]),        // input wire [7 : 0] A_565
  .A_566(A[566]),        // input wire [7 : 0] A_566
  .A_567(A[567]),        // input wire [7 : 0] A_567
  .A_568(A[568]),        // input wire [7 : 0] A_568
  .A_569(A[569]),        // input wire [7 : 0] A_569
  .A_570(A[570]),        // input wire [7 : 0] A_570
  .A_571(A[571]),        // input wire [7 : 0] A_571
  .A_572(A[572]),        // input wire [7 : 0] A_572
  .A_573(A[573]),        // input wire [7 : 0] A_573
  .A_574(A[574]),        // input wire [7 : 0] A_574
  .A_575(A[575]),        // input wire [7 : 0] A_575
  .A_576(A[576]),        // input wire [7 : 0] A_576
  .A_577(A[577]),        // input wire [7 : 0] A_577
  .A_578(A[578]),        // input wire [7 : 0] A_578
  .A_579(A[579]),        // input wire [7 : 0] A_579
  .A_580(A[580]),        // input wire [7 : 0] A_580
  .A_581(A[581]),        // input wire [7 : 0] A_581
  .A_582(A[582]),        // input wire [7 : 0] A_582
  .A_583(A[583]),        // input wire [7 : 0] A_583
  .A_584(A[584]),        // input wire [7 : 0] A_584
  .A_585(A[585]),        // input wire [7 : 0] A_585
  .A_586(A[586]),        // input wire [7 : 0] A_586
  .A_587(A[587]),        // input wire [7 : 0] A_587
  .A_588(A[588]),        // input wire [7 : 0] A_588
  .A_589(A[589]),        // input wire [7 : 0] A_589
  .A_590(A[590]),        // input wire [7 : 0] A_590
  .A_591(A[591]),        // input wire [7 : 0] A_591
  .A_592(A[592]),        // input wire [7 : 0] A_592
  .A_593(A[593]),        // input wire [7 : 0] A_593
  .A_594(A[594]),        // input wire [7 : 0] A_594
  .A_595(A[595]),        // input wire [7 : 0] A_595
  .A_596(A[596]),        // input wire [7 : 0] A_596
  .A_597(A[597]),        // input wire [7 : 0] A_597
  .A_598(A[598]),        // input wire [7 : 0] A_598
  .A_599(A[599]),        // input wire [7 : 0] A_599
  .A_600(A[600]),        // input wire [7 : 0] A_600
  .A_601(A[601]),        // input wire [7 : 0] A_601
  .A_602(A[602]),        // input wire [7 : 0] A_602
  .A_603(A[603]),        // input wire [7 : 0] A_603
  .A_604(A[604]),        // input wire [7 : 0] A_604
  .A_605(A[605]),        // input wire [7 : 0] A_605
  .A_606(A[606]),        // input wire [7 : 0] A_606
  .A_607(A[607]),        // input wire [7 : 0] A_607
  .A_608(A[608]),        // input wire [7 : 0] A_608
  .A_609(A[609]),        // input wire [7 : 0] A_609
  .A_610(A[610]),        // input wire [7 : 0] A_610
  .A_611(A[611]),        // input wire [7 : 0] A_611
  .A_612(A[612]),        // input wire [7 : 0] A_612
  .A_613(A[613]),        // input wire [7 : 0] A_613
  .A_614(A[614]),        // input wire [7 : 0] A_614
  .A_615(A[615]),        // input wire [7 : 0] A_615
  .A_616(A[616]),        // input wire [7 : 0] A_616
  .A_617(A[617]),        // input wire [7 : 0] A_617
  .A_618(A[618]),        // input wire [7 : 0] A_618
  .A_619(A[619]),        // input wire [7 : 0] A_619
  .A_620(A[620]),        // input wire [7 : 0] A_620
  .A_621(A[621]),        // input wire [7 : 0] A_621
  .A_622(A[622]),        // input wire [7 : 0] A_622
  .A_623(A[623]),        // input wire [7 : 0] A_623
  .A_624(A[624]),        // input wire [7 : 0] A_624
  .A_625(A[625]),        // input wire [7 : 0] A_625
  .A_626(A[626]),        // input wire [7 : 0] A_626
  .A_627(A[627]),        // input wire [7 : 0] A_627
  .A_628(A[628]),        // input wire [7 : 0] A_628
  .A_629(A[629]),        // input wire [7 : 0] A_629
  .A_630(A[630]),        // input wire [7 : 0] A_630
  .A_631(A[631]),        // input wire [7 : 0] A_631
  .A_632(A[632]),        // input wire [7 : 0] A_632
  .A_633(A[633]),        // input wire [7 : 0] A_633
  .A_634(A[634]),        // input wire [7 : 0] A_634
  .A_635(A[635]),        // input wire [7 : 0] A_635
  .A_636(A[636]),        // input wire [7 : 0] A_636
  .A_637(A[637]),        // input wire [7 : 0] A_637
  .A_638(A[638]),        // input wire [7 : 0] A_638
  .A_639(A[639]),        // input wire [7 : 0] A_639
  .A_640(A[640]),        // input wire [7 : 0] A_640
  .A_641(A[641]),        // input wire [7 : 0] A_641
  .A_642(A[642]),        // input wire [7 : 0] A_642
  .A_643(A[643]),        // input wire [7 : 0] A_643
  .A_644(A[644]),        // input wire [7 : 0] A_644
  .A_645(A[645]),        // input wire [7 : 0] A_645
  .A_646(A[646]),        // input wire [7 : 0] A_646
  .A_647(A[647]),        // input wire [7 : 0] A_647
  .A_648(A[648]),        // input wire [7 : 0] A_648
  .A_649(A[649]),        // input wire [7 : 0] A_649
  .A_650(A[650]),        // input wire [7 : 0] A_650
  .A_651(A[651]),        // input wire [7 : 0] A_651
  .A_652(A[652]),        // input wire [7 : 0] A_652
  .A_653(A[653]),        // input wire [7 : 0] A_653
  .A_654(A[654]),        // input wire [7 : 0] A_654
  .A_655(A[655]),        // input wire [7 : 0] A_655
  .A_656(A[656]),        // input wire [7 : 0] A_656
  .A_657(A[657]),        // input wire [7 : 0] A_657
  .A_658(A[658]),        // input wire [7 : 0] A_658
  .A_659(A[659]),        // input wire [7 : 0] A_659
  .A_660(A[660]),        // input wire [7 : 0] A_660
  .A_661(A[661]),        // input wire [7 : 0] A_661
  .A_662(A[662]),        // input wire [7 : 0] A_662
  .A_663(A[663]),        // input wire [7 : 0] A_663
  .A_664(A[664]),        // input wire [7 : 0] A_664
  .A_665(A[665]),        // input wire [7 : 0] A_665
  .A_666(A[666]),        // input wire [7 : 0] A_666
  .A_667(A[667]),        // input wire [7 : 0] A_667
  .A_668(A[668]),        // input wire [7 : 0] A_668
  .A_669(A[669]),        // input wire [7 : 0] A_669
  .A_670(A[670]),        // input wire [7 : 0] A_670
  .A_671(A[671]),        // input wire [7 : 0] A_671
  .A_672(A[672]),        // input wire [7 : 0] A_672
  .A_673(A[673]),        // input wire [7 : 0] A_673
  .A_674(A[674]),        // input wire [7 : 0] A_674
  .A_675(A[675]),        // input wire [7 : 0] A_675
  .A_676(A[676]),        // input wire [7 : 0] A_676
  .A_677(A[677]),        // input wire [7 : 0] A_677
  .A_678(A[678]),        // input wire [7 : 0] A_678
  .A_679(A[679]),        // input wire [7 : 0] A_679
  .A_680(A[680]),        // input wire [7 : 0] A_680
  .A_681(A[681]),        // input wire [7 : 0] A_681
  .A_682(A[682]),        // input wire [7 : 0] A_682
  .A_683(A[683]),        // input wire [7 : 0] A_683
  .A_684(A[684]),        // input wire [7 : 0] A_684
  .A_685(A[685]),        // input wire [7 : 0] A_685
  .A_686(A[686]),        // input wire [7 : 0] A_686
  .A_687(A[687]),        // input wire [7 : 0] A_687
  .A_688(A[688]),        // input wire [7 : 0] A_688
  .A_689(A[689]),        // input wire [7 : 0] A_689
  .A_690(A[690]),        // input wire [7 : 0] A_690
  .A_691(A[691]),        // input wire [7 : 0] A_691
  .A_692(A[692]),        // input wire [7 : 0] A_692
  .A_693(A[693]),        // input wire [7 : 0] A_693
  .A_694(A[694]),        // input wire [7 : 0] A_694
  .A_695(A[695]),        // input wire [7 : 0] A_695
  .A_696(A[696]),        // input wire [7 : 0] A_696
  .A_697(A[697]),        // input wire [7 : 0] A_697
  .A_698(A[698]),        // input wire [7 : 0] A_698
  .A_699(A[699]),        // input wire [7 : 0] A_699
  .A_700(A[700]),        // input wire [7 : 0] A_700
  .A_701(A[701]),        // input wire [7 : 0] A_701
  .A_702(A[702]),        // input wire [7 : 0] A_702
  .A_703(A[703]),        // input wire [7 : 0] A_703
  .A_704(A[704]),        // input wire [7 : 0] A_704
  .A_705(A[705]),        // input wire [7 : 0] A_705
  .A_706(A[706]),        // input wire [7 : 0] A_706
  .A_707(A[707]),        // input wire [7 : 0] A_707
  .A_708(A[708]),        // input wire [7 : 0] A_708
  .A_709(A[709]),        // input wire [7 : 0] A_709
  .A_710(A[710]),        // input wire [7 : 0] A_710
  .A_711(A[711]),        // input wire [7 : 0] A_711
  .A_712(A[712]),        // input wire [7 : 0] A_712
  .A_713(A[713]),        // input wire [7 : 0] A_713
  .A_714(A[714]),        // input wire [7 : 0] A_714
  .A_715(A[715]),        // input wire [7 : 0] A_715
  .A_716(A[716]),        // input wire [7 : 0] A_716
  .A_717(A[717]),        // input wire [7 : 0] A_717
  .A_718(A[718]),        // input wire [7 : 0] A_718
  .A_719(A[719]),        // input wire [7 : 0] A_719
  .A_720(A[720]),        // input wire [7 : 0] A_720
  .A_721(A[721]),        // input wire [7 : 0] A_721
  .A_722(A[722]),        // input wire [7 : 0] A_722
  .A_723(A[723]),        // input wire [7 : 0] A_723
  .A_724(A[724]),        // input wire [7 : 0] A_724
  .A_725(A[725]),        // input wire [7 : 0] A_725
  .A_726(A[726]),        // input wire [7 : 0] A_726
  .A_727(A[727]),        // input wire [7 : 0] A_727
  .A_728(A[728]),        // input wire [7 : 0] A_728
  .A_729(A[729]),        // input wire [7 : 0] A_729
  .A_730(A[730]),        // input wire [7 : 0] A_730
  .A_731(A[731]),        // input wire [7 : 0] A_731
  .A_732(A[732]),        // input wire [7 : 0] A_732
  .A_733(A[733]),        // input wire [7 : 0] A_733
  .A_734(A[734]),        // input wire [7 : 0] A_734
  .A_735(A[735]),        // input wire [7 : 0] A_735
  .A_736(A[736]),        // input wire [7 : 0] A_736
  .A_737(A[737]),        // input wire [7 : 0] A_737
  .A_738(A[738]),        // input wire [7 : 0] A_738
  .A_739(A[739]),        // input wire [7 : 0] A_739
  .A_740(A[740]),        // input wire [7 : 0] A_740
  .A_741(A[741]),        // input wire [7 : 0] A_741
  .A_742(A[742]),        // input wire [7 : 0] A_742
  .A_743(A[743]),        // input wire [7 : 0] A_743
  .A_744(A[744]),        // input wire [7 : 0] A_744
  .A_745(A[745]),        // input wire [7 : 0] A_745
  .A_746(A[746]),        // input wire [7 : 0] A_746
  .A_747(A[747]),        // input wire [7 : 0] A_747
  .A_748(A[748]),        // input wire [7 : 0] A_748
  .A_749(A[749]),        // input wire [7 : 0] A_749
  .A_750(A[750]),        // input wire [7 : 0] A_750
  .A_751(A[751]),        // input wire [7 : 0] A_751
  .A_752(A[752]),        // input wire [7 : 0] A_752
  .A_753(A[753]),        // input wire [7 : 0] A_753
  .A_754(A[754]),        // input wire [7 : 0] A_754
  .A_755(A[755]),        // input wire [7 : 0] A_755
  .A_756(A[756]),        // input wire [7 : 0] A_756
  .A_757(A[757]),        // input wire [7 : 0] A_757
  .A_758(A[758]),        // input wire [7 : 0] A_758
  .A_759(A[759]),        // input wire [7 : 0] A_759
  .A_760(A[760]),        // input wire [7 : 0] A_760
  .A_761(A[761]),        // input wire [7 : 0] A_761
  .A_762(A[762]),        // input wire [7 : 0] A_762
  .A_763(A[763]),        // input wire [7 : 0] A_763
  .A_764(A[764]),        // input wire [7 : 0] A_764
  .A_765(A[765]),        // input wire [7 : 0] A_765
  .A_766(A[766]),        // input wire [7 : 0] A_766
  .A_767(A[767]),        // input wire [7 : 0] A_767
  .A_768(A[768]),        // input wire [7 : 0] A_768
  .A_769(A[769]),        // input wire [7 : 0] A_769
  .A_770(A[770]),        // input wire [7 : 0] A_770
  .A_771(A[771]),        // input wire [7 : 0] A_771
  .A_772(A[772]),        // input wire [7 : 0] A_772
  .A_773(A[773]),        // input wire [7 : 0] A_773
  .A_774(A[774]),        // input wire [7 : 0] A_774
  .A_775(A[775]),        // input wire [7 : 0] A_775
  .A_776(A[776]),        // input wire [7 : 0] A_776
  .A_777(A[777]),        // input wire [7 : 0] A_777
  .A_778(A[778]),        // input wire [7 : 0] A_778
  .A_779(A[779]),        // input wire [7 : 0] A_779
  .A_780(A[780]),        // input wire [7 : 0] A_780
  .A_781(A[781]),        // input wire [7 : 0] A_781
  .A_782(A[782]),        // input wire [7 : 0] A_782
  .A_783(A[783]),        // input wire [7 : 0] A_783
  .A_784(A[784]),        // input wire [7 : 0] A_784
  .A_785(A[785]),        // input wire [7 : 0] A_785
  .A_786(A[786]),        // input wire [7 : 0] A_786
  .A_787(A[787]),        // input wire [7 : 0] A_787
  .A_788(A[788]),        // input wire [7 : 0] A_788
  .A_789(A[789]),        // input wire [7 : 0] A_789
  .A_790(A[790]),        // input wire [7 : 0] A_790
  .A_791(A[791]),        // input wire [7 : 0] A_791
  .A_792(A[792]),        // input wire [7 : 0] A_792
  .A_793(A[793]),        // input wire [7 : 0] A_793
  .A_794(A[794]),        // input wire [7 : 0] A_794
  .A_795(A[795]),        // input wire [7 : 0] A_795
  .A_796(A[796]),        // input wire [7 : 0] A_796
  .A_797(A[797]),        // input wire [7 : 0] A_797
  .A_798(A[798]),        // input wire [7 : 0] A_798
  .A_799(A[799]),        // input wire [7 : 0] A_799
  .A_800(A[800]),        // input wire [7 : 0] A_800
  .A_801(A[801]),        // input wire [7 : 0] A_801
  .A_802(A[802]),        // input wire [7 : 0] A_802
  .A_803(A[803]),        // input wire [7 : 0] A_803
  .A_804(A[804]),        // input wire [7 : 0] A_804
  .A_805(A[805]),        // input wire [7 : 0] A_805
  .A_806(A[806]),        // input wire [7 : 0] A_806
  .A_807(A[807]),        // input wire [7 : 0] A_807
  .A_808(A[808]),        // input wire [7 : 0] A_808
  .A_809(A[809]),        // input wire [7 : 0] A_809
  .A_810(A[810]),        // input wire [7 : 0] A_810
  .A_811(A[811]),        // input wire [7 : 0] A_811
  .A_812(A[812]),        // input wire [7 : 0] A_812
  .A_813(A[813]),        // input wire [7 : 0] A_813
  .A_814(A[814]),        // input wire [7 : 0] A_814
  .A_815(A[815]),        // input wire [7 : 0] A_815
  .A_816(A[816]),        // input wire [7 : 0] A_816
  .A_817(A[817]),        // input wire [7 : 0] A_817
  .A_818(A[818]),        // input wire [7 : 0] A_818
  .A_819(A[819]),        // input wire [7 : 0] A_819
  .A_820(A[820]),        // input wire [7 : 0] A_820
  .A_821(A[821]),        // input wire [7 : 0] A_821
  .A_822(A[822]),        // input wire [7 : 0] A_822
  .A_823(A[823]),        // input wire [7 : 0] A_823
  .A_824(A[824]),        // input wire [7 : 0] A_824
  .A_825(A[825]),        // input wire [7 : 0] A_825
  .A_826(A[826]),        // input wire [7 : 0] A_826
  .A_827(A[827]),        // input wire [7 : 0] A_827
  .A_828(A[828]),        // input wire [7 : 0] A_828
  .A_829(A[829]),        // input wire [7 : 0] A_829
  .A_830(A[830]),        // input wire [7 : 0] A_830
  .A_831(A[831]),        // input wire [7 : 0] A_831
  .A_832(A[832]),        // input wire [7 : 0] A_832
  .A_833(A[833]),        // input wire [7 : 0] A_833
  .A_834(A[834]),        // input wire [7 : 0] A_834
  .A_835(A[835]),        // input wire [7 : 0] A_835
  .A_836(A[836]),        // input wire [7 : 0] A_836
  .A_837(A[837]),        // input wire [7 : 0] A_837
  .A_838(A[838]),        // input wire [7 : 0] A_838
  .A_839(A[839]),        // input wire [7 : 0] A_839
  .A_840(A[840]),        // input wire [7 : 0] A_840
  .A_841(A[841]),        // input wire [7 : 0] A_841
  .A_842(A[842]),        // input wire [7 : 0] A_842
  .A_843(A[843]),        // input wire [7 : 0] A_843
  .A_844(A[844]),        // input wire [7 : 0] A_844
  .A_845(A[845]),        // input wire [7 : 0] A_845
  .A_846(A[846]),        // input wire [7 : 0] A_846
  .A_847(A[847]),        // input wire [7 : 0] A_847
  .A_848(A[848]),        // input wire [7 : 0] A_848
  .A_849(A[849]),        // input wire [7 : 0] A_849
  .A_850(A[850]),        // input wire [7 : 0] A_850
  .A_851(A[851]),        // input wire [7 : 0] A_851
  .A_852(A[852]),        // input wire [7 : 0] A_852
  .A_853(A[853]),        // input wire [7 : 0] A_853
  .A_854(A[854]),        // input wire [7 : 0] A_854
  .A_855(A[855]),        // input wire [7 : 0] A_855
  .A_856(A[856]),        // input wire [7 : 0] A_856
  .A_857(A[857]),        // input wire [7 : 0] A_857
  .A_858(A[858]),        // input wire [7 : 0] A_858
  .A_859(A[859]),        // input wire [7 : 0] A_859
  .A_860(A[860]),        // input wire [7 : 0] A_860
  .A_861(A[861]),        // input wire [7 : 0] A_861
  .A_862(A[862]),        // input wire [7 : 0] A_862
  .A_863(A[863]),        // input wire [7 : 0] A_863
  .A_864(A[864]),        // input wire [7 : 0] A_864
  .A_865(A[865]),        // input wire [7 : 0] A_865
  .A_866(A[866]),        // input wire [7 : 0] A_866
  .A_867(A[867]),        // input wire [7 : 0] A_867
  .A_868(A[868]),        // input wire [7 : 0] A_868
  .A_869(A[869]),        // input wire [7 : 0] A_869
  .A_870(A[870]),        // input wire [7 : 0] A_870
  .A_871(A[871]),        // input wire [7 : 0] A_871
  .A_872(A[872]),        // input wire [7 : 0] A_872
  .A_873(A[873]),        // input wire [7 : 0] A_873
  .A_874(A[874]),        // input wire [7 : 0] A_874
  .A_875(A[875]),        // input wire [7 : 0] A_875
  .A_876(A[876]),        // input wire [7 : 0] A_876
  .A_877(A[877]),        // input wire [7 : 0] A_877
  .A_878(A[878]),        // input wire [7 : 0] A_878
  .A_879(A[879]),        // input wire [7 : 0] A_879
  .A_880(A[880]),        // input wire [7 : 0] A_880
  .A_881(A[881]),        // input wire [7 : 0] A_881
  .A_882(A[882]),        // input wire [7 : 0] A_882
  .A_883(A[883]),        // input wire [7 : 0] A_883
  .A_884(A[884]),        // input wire [7 : 0] A_884
  .A_885(A[885]),        // input wire [7 : 0] A_885
  .A_886(A[886]),        // input wire [7 : 0] A_886
  .A_887(A[887]),        // input wire [7 : 0] A_887
  .A_888(A[888]),        // input wire [7 : 0] A_888
  .A_889(A[889]),        // input wire [7 : 0] A_889
  .A_890(A[890]),        // input wire [7 : 0] A_890
  .A_891(A[891]),        // input wire [7 : 0] A_891
  .A_892(A[892]),        // input wire [7 : 0] A_892
  .A_893(A[893]),        // input wire [7 : 0] A_893
  .A_894(A[894]),        // input wire [7 : 0] A_894
  .A_895(A[895]),        // input wire [7 : 0] A_895
  .A_896(A[896]),        // input wire [7 : 0] A_896
  .A_897(A[897]),        // input wire [7 : 0] A_897
  .A_898(A[898]),        // input wire [7 : 0] A_898
  .A_899(A[899]),        // input wire [7 : 0] A_899
  .A_900(A[900]),        // input wire [7 : 0] A_900
  .A_901(A[901]),        // input wire [7 : 0] A_901
  .A_902(A[902]),        // input wire [7 : 0] A_902
  .A_903(A[903]),        // input wire [7 : 0] A_903
  .A_904(A[904]),        // input wire [7 : 0] A_904
  .A_905(A[905]),        // input wire [7 : 0] A_905
  .A_906(A[906]),        // input wire [7 : 0] A_906
  .A_907(A[907]),        // input wire [7 : 0] A_907
  .A_908(A[908]),        // input wire [7 : 0] A_908
  .A_909(A[909]),        // input wire [7 : 0] A_909
  .A_910(A[910]),        // input wire [7 : 0] A_910
  .A_911(A[911]),        // input wire [7 : 0] A_911
  .A_912(A[912]),        // input wire [7 : 0] A_912
  .A_913(A[913]),        // input wire [7 : 0] A_913
  .A_914(A[914]),        // input wire [7 : 0] A_914
  .A_915(A[915]),        // input wire [7 : 0] A_915
  .A_916(A[916]),        // input wire [7 : 0] A_916
  .A_917(A[917]),        // input wire [7 : 0] A_917
  .A_918(A[918]),        // input wire [7 : 0] A_918
  .A_919(A[919]),        // input wire [7 : 0] A_919
  .A_920(A[920]),        // input wire [7 : 0] A_920
  .A_921(A[921]),        // input wire [7 : 0] A_921
  .A_922(A[922]),        // input wire [7 : 0] A_922
  .A_923(A[923]),        // input wire [7 : 0] A_923
  .A_924(A[924]),        // input wire [7 : 0] A_924
  .A_925(A[925]),        // input wire [7 : 0] A_925
  .A_926(A[926]),        // input wire [7 : 0] A_926
  .A_927(A[927]),        // input wire [7 : 0] A_927
  .A_928(A[928]),        // input wire [7 : 0] A_928
  .A_929(A[929]),        // input wire [7 : 0] A_929
  .A_930(A[930]),        // input wire [7 : 0] A_930
  .A_931(A[931]),        // input wire [7 : 0] A_931
  .A_932(A[932]),        // input wire [7 : 0] A_932
  .A_933(A[933]),        // input wire [7 : 0] A_933
  .A_934(A[934]),        // input wire [7 : 0] A_934
  .A_935(A[935]),        // input wire [7 : 0] A_935
  .A_936(A[936]),        // input wire [7 : 0] A_936
  .A_937(A[937]),        // input wire [7 : 0] A_937
  .A_938(A[938]),        // input wire [7 : 0] A_938
  .A_939(A[939]),        // input wire [7 : 0] A_939
  .A_940(A[940]),        // input wire [7 : 0] A_940
  .A_941(A[941]),        // input wire [7 : 0] A_941
  .A_942(A[942]),        // input wire [7 : 0] A_942
  .A_943(A[943]),        // input wire [7 : 0] A_943
  .A_944(A[944]),        // input wire [7 : 0] A_944
  .A_945(A[945]),        // input wire [7 : 0] A_945
  .A_946(A[946]),        // input wire [7 : 0] A_946
  .A_947(A[947]),        // input wire [7 : 0] A_947
  .A_948(A[948]),        // input wire [7 : 0] A_948
  .A_949(A[949]),        // input wire [7 : 0] A_949
  .A_950(A[950]),        // input wire [7 : 0] A_950
  .A_951(A[951]),        // input wire [7 : 0] A_951
  .A_952(A[952]),        // input wire [7 : 0] A_952
  .A_953(A[953]),        // input wire [7 : 0] A_953
  .A_954(A[954]),        // input wire [7 : 0] A_954
  .A_955(A[955]),        // input wire [7 : 0] A_955
  .A_956(A[956]),        // input wire [7 : 0] A_956
  .A_957(A[957]),        // input wire [7 : 0] A_957
  .A_958(A[958]),        // input wire [7 : 0] A_958
  .A_959(A[959]),        // input wire [7 : 0] A_959
  .A_960(A[960]),        // input wire [7 : 0] A_960
  .A_961(A[961]),        // input wire [7 : 0] A_961
  .A_962(A[962]),        // input wire [7 : 0] A_962
  .A_963(A[963]),        // input wire [7 : 0] A_963
  .A_964(A[964]),        // input wire [7 : 0] A_964
  .A_965(A[965]),        // input wire [7 : 0] A_965
  .A_966(A[966]),        // input wire [7 : 0] A_966
  .A_967(A[967]),        // input wire [7 : 0] A_967
  .A_968(A[968]),        // input wire [7 : 0] A_968
  .A_969(A[969]),        // input wire [7 : 0] A_969
  .A_970(A[970]),        // input wire [7 : 0] A_970
  .A_971(A[971]),        // input wire [7 : 0] A_971
  .A_972(A[972]),        // input wire [7 : 0] A_972
  .A_973(A[973]),        // input wire [7 : 0] A_973
  .A_974(A[974]),        // input wire [7 : 0] A_974
  .A_975(A[975]),        // input wire [7 : 0] A_975
  .A_976(A[976]),        // input wire [7 : 0] A_976
  .A_977(A[977]),        // input wire [7 : 0] A_977
  .A_978(A[978]),        // input wire [7 : 0] A_978
  .A_979(A[979]),        // input wire [7 : 0] A_979
  .A_980(A[980]),        // input wire [7 : 0] A_980
  .A_981(A[981]),        // input wire [7 : 0] A_981
  .A_982(A[982]),        // input wire [7 : 0] A_982
  .A_983(A[983]),        // input wire [7 : 0] A_983
  .A_984(A[984]),        // input wire [7 : 0] A_984
  .A_985(A[985]),        // input wire [7 : 0] A_985
  .A_986(A[986]),        // input wire [7 : 0] A_986
  .A_987(A[987]),        // input wire [7 : 0] A_987
  .A_988(A[988]),        // input wire [7 : 0] A_988
  .A_989(A[989]),        // input wire [7 : 0] A_989
  .A_990(A[990]),        // input wire [7 : 0] A_990
  .A_991(A[991]),        // input wire [7 : 0] A_991
  .A_992(A[992]),        // input wire [7 : 0] A_992
  .A_993(A[993]),        // input wire [7 : 0] A_993
  .A_994(A[994]),        // input wire [7 : 0] A_994
  .A_995(A[995]),        // input wire [7 : 0] A_995
  .A_996(A[996]),        // input wire [7 : 0] A_996
  .A_997(A[997]),        // input wire [7 : 0] A_997
  .A_998(A[998]),        // input wire [7 : 0] A_998
  .A_999(A[999]),        // input wire [7 : 0] A_999
  .A_1000(A[1000]),      // input wire [7 : 0] A_1000
  .A_1001(A[1001]),      // input wire [7 : 0] A_1001
  .A_1002(A[1002]),      // input wire [7 : 0] A_1002
  .A_1003(A[1003]),      // input wire [7 : 0] A_1003
  .A_1004(A[1004]),      // input wire [7 : 0] A_1004
  .A_1005(A[1005]),      // input wire [7 : 0] A_1005
  .A_1006(A[1006]),      // input wire [7 : 0] A_1006
  .A_1007(A[1007]),      // input wire [7 : 0] A_1007
  .A_1008(A[1008]),      // input wire [7 : 0] A_1008
  .A_1009(A[1009]),      // input wire [7 : 0] A_1009
  .A_1010(A[1010]),      // input wire [7 : 0] A_1010
  .A_1011(A[1011]),      // input wire [7 : 0] A_1011
  .A_1012(A[1012]),      // input wire [7 : 0] A_1012
  .A_1013(A[1013]),      // input wire [7 : 0] A_1013
  .A_1014(A[1014]),      // input wire [7 : 0] A_1014
  .A_1015(A[1015]),      // input wire [7 : 0] A_1015
  .A_1016(A[1016]),      // input wire [7 : 0] A_1016
  .A_1017(A[1017]),      // input wire [7 : 0] A_1017
  .A_1018(A[1018]),      // input wire [7 : 0] A_1018
  .A_1019(A[1019]),      // input wire [7 : 0] A_1019
  .A_1020(A[1020]),      // input wire [7 : 0] A_1020
  .A_1021(A[1021]),      // input wire [7 : 0] A_1021
  .A_1022(A[1022]),      // input wire [7 : 0] A_1022
  .A_1023(A[1023]),      // input wire [7 : 0] A_1023
  .B_0(B[0]),            // input wire [7 : 0] B_0
  .B_1(B[1]),            // input wire [7 : 0] B_1
  .B_2(B[2]),            // input wire [7 : 0] B_2
  .B_3(B[3]),            // input wire [7 : 0] B_3
  .B_4(B[4]),            // input wire [7 : 0] B_4
  .B_5(B[5]),            // input wire [7 : 0] B_5
  .B_6(B[6]),            // input wire [7 : 0] B_6
  .B_7(B[7]),            // input wire [7 : 0] B_7
  .B_8(B[8]),            // input wire [7 : 0] B_8
  .B_9(B[9]),            // input wire [7 : 0] B_9
  .B_10(B[10]),          // input wire [7 : 0] B_10
  .B_11(B[11]),          // input wire [7 : 0] B_11
  .B_12(B[12]),          // input wire [7 : 0] B_12
  .B_13(B[13]),          // input wire [7 : 0] B_13
  .B_14(B[14]),          // input wire [7 : 0] B_14
  .B_15(B[15]),          // input wire [7 : 0] B_15
  .B_16(B[16]),          // input wire [7 : 0] B_16
  .B_17(B[17]),          // input wire [7 : 0] B_17
  .B_18(B[18]),          // input wire [7 : 0] B_18
  .B_19(B[19]),          // input wire [7 : 0] B_19
  .B_20(B[20]),          // input wire [7 : 0] B_20
  .B_21(B[21]),          // input wire [7 : 0] B_21
  .B_22(B[22]),          // input wire [7 : 0] B_22
  .B_23(B[23]),          // input wire [7 : 0] B_23
  .B_24(B[24]),          // input wire [7 : 0] B_24
  .B_25(B[25]),          // input wire [7 : 0] B_25
  .B_26(B[26]),          // input wire [7 : 0] B_26
  .B_27(B[27]),          // input wire [7 : 0] B_27
  .B_28(B[28]),          // input wire [7 : 0] B_28
  .B_29(B[29]),          // input wire [7 : 0] B_29
  .B_30(B[30]),          // input wire [7 : 0] B_30
  .B_31(B[31]),          // input wire [7 : 0] B_31
  .B_32(B[32]),          // input wire [7 : 0] B_32
  .B_33(B[33]),          // input wire [7 : 0] B_33
  .B_34(B[34]),          // input wire [7 : 0] B_34
  .B_35(B[35]),          // input wire [7 : 0] B_35
  .B_36(B[36]),          // input wire [7 : 0] B_36
  .B_37(B[37]),          // input wire [7 : 0] B_37
  .B_38(B[38]),          // input wire [7 : 0] B_38
  .B_39(B[39]),          // input wire [7 : 0] B_39
  .B_40(B[40]),          // input wire [7 : 0] B_40
  .B_41(B[41]),          // input wire [7 : 0] B_41
  .B_42(B[42]),          // input wire [7 : 0] B_42
  .B_43(B[43]),          // input wire [7 : 0] B_43
  .B_44(B[44]),          // input wire [7 : 0] B_44
  .B_45(B[45]),          // input wire [7 : 0] B_45
  .B_46(B[46]),          // input wire [7 : 0] B_46
  .B_47(B[47]),          // input wire [7 : 0] B_47
  .B_48(B[48]),          // input wire [7 : 0] B_48
  .B_49(B[49]),          // input wire [7 : 0] B_49
  .B_50(B[50]),          // input wire [7 : 0] B_50
  .B_51(B[51]),          // input wire [7 : 0] B_51
  .B_52(B[52]),          // input wire [7 : 0] B_52
  .B_53(B[53]),          // input wire [7 : 0] B_53
  .B_54(B[54]),          // input wire [7 : 0] B_54
  .B_55(B[55]),          // input wire [7 : 0] B_55
  .B_56(B[56]),          // input wire [7 : 0] B_56
  .B_57(B[57]),          // input wire [7 : 0] B_57
  .B_58(B[58]),          // input wire [7 : 0] B_58
  .B_59(B[59]),          // input wire [7 : 0] B_59
  .B_60(B[60]),          // input wire [7 : 0] B_60
  .B_61(B[61]),          // input wire [7 : 0] B_61
  .B_62(B[62]),          // input wire [7 : 0] B_62
  .B_63(B[63]),          // input wire [7 : 0] B_63
  .B_64(B[64]),          // input wire [7 : 0] B_64
  .B_65(B[65]),          // input wire [7 : 0] B_65
  .B_66(B[66]),          // input wire [7 : 0] B_66
  .B_67(B[67]),          // input wire [7 : 0] B_67
  .B_68(B[68]),          // input wire [7 : 0] B_68
  .B_69(B[69]),          // input wire [7 : 0] B_69
  .B_70(B[70]),          // input wire [7 : 0] B_70
  .B_71(B[71]),          // input wire [7 : 0] B_71
  .B_72(B[72]),          // input wire [7 : 0] B_72
  .B_73(B[73]),          // input wire [7 : 0] B_73
  .B_74(B[74]),          // input wire [7 : 0] B_74
  .B_75(B[75]),          // input wire [7 : 0] B_75
  .B_76(B[76]),          // input wire [7 : 0] B_76
  .B_77(B[77]),          // input wire [7 : 0] B_77
  .B_78(B[78]),          // input wire [7 : 0] B_78
  .B_79(B[79]),          // input wire [7 : 0] B_79
  .B_80(B[80]),          // input wire [7 : 0] B_80
  .B_81(B[81]),          // input wire [7 : 0] B_81
  .B_82(B[82]),          // input wire [7 : 0] B_82
  .B_83(B[83]),          // input wire [7 : 0] B_83
  .B_84(B[84]),          // input wire [7 : 0] B_84
  .B_85(B[85]),          // input wire [7 : 0] B_85
  .B_86(B[86]),          // input wire [7 : 0] B_86
  .B_87(B[87]),          // input wire [7 : 0] B_87
  .B_88(B[88]),          // input wire [7 : 0] B_88
  .B_89(B[89]),          // input wire [7 : 0] B_89
  .B_90(B[90]),          // input wire [7 : 0] B_90
  .B_91(B[91]),          // input wire [7 : 0] B_91
  .B_92(B[92]),          // input wire [7 : 0] B_92
  .B_93(B[93]),          // input wire [7 : 0] B_93
  .B_94(B[94]),          // input wire [7 : 0] B_94
  .B_95(B[95]),          // input wire [7 : 0] B_95
  .B_96(B[96]),          // input wire [7 : 0] B_96
  .B_97(B[97]),          // input wire [7 : 0] B_97
  .B_98(B[98]),          // input wire [7 : 0] B_98
  .B_99(B[99]),          // input wire [7 : 0] B_99
  .B_100(B[100]),        // input wire [7 : 0] B_100
  .B_101(B[101]),        // input wire [7 : 0] B_101
  .B_102(B[102]),        // input wire [7 : 0] B_102
  .B_103(B[103]),        // input wire [7 : 0] B_103
  .B_104(B[104]),        // input wire [7 : 0] B_104
  .B_105(B[105]),        // input wire [7 : 0] B_105
  .B_106(B[106]),        // input wire [7 : 0] B_106
  .B_107(B[107]),        // input wire [7 : 0] B_107
  .B_108(B[108]),        // input wire [7 : 0] B_108
  .B_109(B[109]),        // input wire [7 : 0] B_109
  .B_110(B[110]),        // input wire [7 : 0] B_110
  .B_111(B[111]),        // input wire [7 : 0] B_111
  .B_112(B[112]),        // input wire [7 : 0] B_112
  .B_113(B[113]),        // input wire [7 : 0] B_113
  .B_114(B[114]),        // input wire [7 : 0] B_114
  .B_115(B[115]),        // input wire [7 : 0] B_115
  .B_116(B[116]),        // input wire [7 : 0] B_116
  .B_117(B[117]),        // input wire [7 : 0] B_117
  .B_118(B[118]),        // input wire [7 : 0] B_118
  .B_119(B[119]),        // input wire [7 : 0] B_119
  .B_120(B[120]),        // input wire [7 : 0] B_120
  .B_121(B[121]),        // input wire [7 : 0] B_121
  .B_122(B[122]),        // input wire [7 : 0] B_122
  .B_123(B[123]),        // input wire [7 : 0] B_123
  .B_124(B[124]),        // input wire [7 : 0] B_124
  .B_125(B[125]),        // input wire [7 : 0] B_125
  .B_126(B[126]),        // input wire [7 : 0] B_126
  .B_127(B[127]),        // input wire [7 : 0] B_127
  .B_128(B[128]),        // input wire [7 : 0] B_128
  .B_129(B[129]),        // input wire [7 : 0] B_129
  .B_130(B[130]),        // input wire [7 : 0] B_130
  .B_131(B[131]),        // input wire [7 : 0] B_131
  .B_132(B[132]),        // input wire [7 : 0] B_132
  .B_133(B[133]),        // input wire [7 : 0] B_133
  .B_134(B[134]),        // input wire [7 : 0] B_134
  .B_135(B[135]),        // input wire [7 : 0] B_135
  .B_136(B[136]),        // input wire [7 : 0] B_136
  .B_137(B[137]),        // input wire [7 : 0] B_137
  .B_138(B[138]),        // input wire [7 : 0] B_138
  .B_139(B[139]),        // input wire [7 : 0] B_139
  .B_140(B[140]),        // input wire [7 : 0] B_140
  .B_141(B[141]),        // input wire [7 : 0] B_141
  .B_142(B[142]),        // input wire [7 : 0] B_142
  .B_143(B[143]),        // input wire [7 : 0] B_143
  .B_144(B[144]),        // input wire [7 : 0] B_144
  .B_145(B[145]),        // input wire [7 : 0] B_145
  .B_146(B[146]),        // input wire [7 : 0] B_146
  .B_147(B[147]),        // input wire [7 : 0] B_147
  .B_148(B[148]),        // input wire [7 : 0] B_148
  .B_149(B[149]),        // input wire [7 : 0] B_149
  .B_150(B[150]),        // input wire [7 : 0] B_150
  .B_151(B[151]),        // input wire [7 : 0] B_151
  .B_152(B[152]),        // input wire [7 : 0] B_152
  .B_153(B[153]),        // input wire [7 : 0] B_153
  .B_154(B[154]),        // input wire [7 : 0] B_154
  .B_155(B[155]),        // input wire [7 : 0] B_155
  .B_156(B[156]),        // input wire [7 : 0] B_156
  .B_157(B[157]),        // input wire [7 : 0] B_157
  .B_158(B[158]),        // input wire [7 : 0] B_158
  .B_159(B[159]),        // input wire [7 : 0] B_159
  .B_160(B[160]),        // input wire [7 : 0] B_160
  .B_161(B[161]),        // input wire [7 : 0] B_161
  .B_162(B[162]),        // input wire [7 : 0] B_162
  .B_163(B[163]),        // input wire [7 : 0] B_163
  .B_164(B[164]),        // input wire [7 : 0] B_164
  .B_165(B[165]),        // input wire [7 : 0] B_165
  .B_166(B[166]),        // input wire [7 : 0] B_166
  .B_167(B[167]),        // input wire [7 : 0] B_167
  .B_168(B[168]),        // input wire [7 : 0] B_168
  .B_169(B[169]),        // input wire [7 : 0] B_169
  .B_170(B[170]),        // input wire [7 : 0] B_170
  .B_171(B[171]),        // input wire [7 : 0] B_171
  .B_172(B[172]),        // input wire [7 : 0] B_172
  .B_173(B[173]),        // input wire [7 : 0] B_173
  .B_174(B[174]),        // input wire [7 : 0] B_174
  .B_175(B[175]),        // input wire [7 : 0] B_175
  .B_176(B[176]),        // input wire [7 : 0] B_176
  .B_177(B[177]),        // input wire [7 : 0] B_177
  .B_178(B[178]),        // input wire [7 : 0] B_178
  .B_179(B[179]),        // input wire [7 : 0] B_179
  .B_180(B[180]),        // input wire [7 : 0] B_180
  .B_181(B[181]),        // input wire [7 : 0] B_181
  .B_182(B[182]),        // input wire [7 : 0] B_182
  .B_183(B[183]),        // input wire [7 : 0] B_183
  .B_184(B[184]),        // input wire [7 : 0] B_184
  .B_185(B[185]),        // input wire [7 : 0] B_185
  .B_186(B[186]),        // input wire [7 : 0] B_186
  .B_187(B[187]),        // input wire [7 : 0] B_187
  .B_188(B[188]),        // input wire [7 : 0] B_188
  .B_189(B[189]),        // input wire [7 : 0] B_189
  .B_190(B[190]),        // input wire [7 : 0] B_190
  .B_191(B[191]),        // input wire [7 : 0] B_191
  .B_192(B[192]),        // input wire [7 : 0] B_192
  .B_193(B[193]),        // input wire [7 : 0] B_193
  .B_194(B[194]),        // input wire [7 : 0] B_194
  .B_195(B[195]),        // input wire [7 : 0] B_195
  .B_196(B[196]),        // input wire [7 : 0] B_196
  .B_197(B[197]),        // input wire [7 : 0] B_197
  .B_198(B[198]),        // input wire [7 : 0] B_198
  .B_199(B[199]),        // input wire [7 : 0] B_199
  .B_200(B[200]),        // input wire [7 : 0] B_200
  .B_201(B[201]),        // input wire [7 : 0] B_201
  .B_202(B[202]),        // input wire [7 : 0] B_202
  .B_203(B[203]),        // input wire [7 : 0] B_203
  .B_204(B[204]),        // input wire [7 : 0] B_204
  .B_205(B[205]),        // input wire [7 : 0] B_205
  .B_206(B[206]),        // input wire [7 : 0] B_206
  .B_207(B[207]),        // input wire [7 : 0] B_207
  .B_208(B[208]),        // input wire [7 : 0] B_208
  .B_209(B[209]),        // input wire [7 : 0] B_209
  .B_210(B[210]),        // input wire [7 : 0] B_210
  .B_211(B[211]),        // input wire [7 : 0] B_211
  .B_212(B[212]),        // input wire [7 : 0] B_212
  .B_213(B[213]),        // input wire [7 : 0] B_213
  .B_214(B[214]),        // input wire [7 : 0] B_214
  .B_215(B[215]),        // input wire [7 : 0] B_215
  .B_216(B[216]),        // input wire [7 : 0] B_216
  .B_217(B[217]),        // input wire [7 : 0] B_217
  .B_218(B[218]),        // input wire [7 : 0] B_218
  .B_219(B[219]),        // input wire [7 : 0] B_219
  .B_220(B[220]),        // input wire [7 : 0] B_220
  .B_221(B[221]),        // input wire [7 : 0] B_221
  .B_222(B[222]),        // input wire [7 : 0] B_222
  .B_223(B[223]),        // input wire [7 : 0] B_223
  .B_224(B[224]),        // input wire [7 : 0] B_224
  .B_225(B[225]),        // input wire [7 : 0] B_225
  .B_226(B[226]),        // input wire [7 : 0] B_226
  .B_227(B[227]),        // input wire [7 : 0] B_227
  .B_228(B[228]),        // input wire [7 : 0] B_228
  .B_229(B[229]),        // input wire [7 : 0] B_229
  .B_230(B[230]),        // input wire [7 : 0] B_230
  .B_231(B[231]),        // input wire [7 : 0] B_231
  .B_232(B[232]),        // input wire [7 : 0] B_232
  .B_233(B[233]),        // input wire [7 : 0] B_233
  .B_234(B[234]),        // input wire [7 : 0] B_234
  .B_235(B[235]),        // input wire [7 : 0] B_235
  .B_236(B[236]),        // input wire [7 : 0] B_236
  .B_237(B[237]),        // input wire [7 : 0] B_237
  .B_238(B[238]),        // input wire [7 : 0] B_238
  .B_239(B[239]),        // input wire [7 : 0] B_239
  .B_240(B[240]),        // input wire [7 : 0] B_240
  .B_241(B[241]),        // input wire [7 : 0] B_241
  .B_242(B[242]),        // input wire [7 : 0] B_242
  .B_243(B[243]),        // input wire [7 : 0] B_243
  .B_244(B[244]),        // input wire [7 : 0] B_244
  .B_245(B[245]),        // input wire [7 : 0] B_245
  .B_246(B[246]),        // input wire [7 : 0] B_246
  .B_247(B[247]),        // input wire [7 : 0] B_247
  .B_248(B[248]),        // input wire [7 : 0] B_248
  .B_249(B[249]),        // input wire [7 : 0] B_249
  .B_250(B[250]),        // input wire [7 : 0] B_250
  .B_251(B[251]),        // input wire [7 : 0] B_251
  .B_252(B[252]),        // input wire [7 : 0] B_252
  .B_253(B[253]),        // input wire [7 : 0] B_253
  .B_254(B[254]),        // input wire [7 : 0] B_254
  .B_255(B[255]),        // input wire [7 : 0] B_255
  .B_256(B[256]),        // input wire [7 : 0] B_256
  .B_257(B[257]),        // input wire [7 : 0] B_257
  .B_258(B[258]),        // input wire [7 : 0] B_258
  .B_259(B[259]),        // input wire [7 : 0] B_259
  .B_260(B[260]),        // input wire [7 : 0] B_260
  .B_261(B[261]),        // input wire [7 : 0] B_261
  .B_262(B[262]),        // input wire [7 : 0] B_262
  .B_263(B[263]),        // input wire [7 : 0] B_263
  .B_264(B[264]),        // input wire [7 : 0] B_264
  .B_265(B[265]),        // input wire [7 : 0] B_265
  .B_266(B[266]),        // input wire [7 : 0] B_266
  .B_267(B[267]),        // input wire [7 : 0] B_267
  .B_268(B[268]),        // input wire [7 : 0] B_268
  .B_269(B[269]),        // input wire [7 : 0] B_269
  .B_270(B[270]),        // input wire [7 : 0] B_270
  .B_271(B[271]),        // input wire [7 : 0] B_271
  .B_272(B[272]),        // input wire [7 : 0] B_272
  .B_273(B[273]),        // input wire [7 : 0] B_273
  .B_274(B[274]),        // input wire [7 : 0] B_274
  .B_275(B[275]),        // input wire [7 : 0] B_275
  .B_276(B[276]),        // input wire [7 : 0] B_276
  .B_277(B[277]),        // input wire [7 : 0] B_277
  .B_278(B[278]),        // input wire [7 : 0] B_278
  .B_279(B[279]),        // input wire [7 : 0] B_279
  .B_280(B[280]),        // input wire [7 : 0] B_280
  .B_281(B[281]),        // input wire [7 : 0] B_281
  .B_282(B[282]),        // input wire [7 : 0] B_282
  .B_283(B[283]),        // input wire [7 : 0] B_283
  .B_284(B[284]),        // input wire [7 : 0] B_284
  .B_285(B[285]),        // input wire [7 : 0] B_285
  .B_286(B[286]),        // input wire [7 : 0] B_286
  .B_287(B[287]),        // input wire [7 : 0] B_287
  .B_288(B[288]),        // input wire [7 : 0] B_288
  .B_289(B[289]),        // input wire [7 : 0] B_289
  .B_290(B[290]),        // input wire [7 : 0] B_290
  .B_291(B[291]),        // input wire [7 : 0] B_291
  .B_292(B[292]),        // input wire [7 : 0] B_292
  .B_293(B[293]),        // input wire [7 : 0] B_293
  .B_294(B[294]),        // input wire [7 : 0] B_294
  .B_295(B[295]),        // input wire [7 : 0] B_295
  .B_296(B[296]),        // input wire [7 : 0] B_296
  .B_297(B[297]),        // input wire [7 : 0] B_297
  .B_298(B[298]),        // input wire [7 : 0] B_298
  .B_299(B[299]),        // input wire [7 : 0] B_299
  .B_300(B[300]),        // input wire [7 : 0] B_300
  .B_301(B[301]),        // input wire [7 : 0] B_301
  .B_302(B[302]),        // input wire [7 : 0] B_302
  .B_303(B[303]),        // input wire [7 : 0] B_303
  .B_304(B[304]),        // input wire [7 : 0] B_304
  .B_305(B[305]),        // input wire [7 : 0] B_305
  .B_306(B[306]),        // input wire [7 : 0] B_306
  .B_307(B[307]),        // input wire [7 : 0] B_307
  .B_308(B[308]),        // input wire [7 : 0] B_308
  .B_309(B[309]),        // input wire [7 : 0] B_309
  .B_310(B[310]),        // input wire [7 : 0] B_310
  .B_311(B[311]),        // input wire [7 : 0] B_311
  .B_312(B[312]),        // input wire [7 : 0] B_312
  .B_313(B[313]),        // input wire [7 : 0] B_313
  .B_314(B[314]),        // input wire [7 : 0] B_314
  .B_315(B[315]),        // input wire [7 : 0] B_315
  .B_316(B[316]),        // input wire [7 : 0] B_316
  .B_317(B[317]),        // input wire [7 : 0] B_317
  .B_318(B[318]),        // input wire [7 : 0] B_318
  .B_319(B[319]),        // input wire [7 : 0] B_319
  .B_320(B[320]),        // input wire [7 : 0] B_320
  .B_321(B[321]),        // input wire [7 : 0] B_321
  .B_322(B[322]),        // input wire [7 : 0] B_322
  .B_323(B[323]),        // input wire [7 : 0] B_323
  .B_324(B[324]),        // input wire [7 : 0] B_324
  .B_325(B[325]),        // input wire [7 : 0] B_325
  .B_326(B[326]),        // input wire [7 : 0] B_326
  .B_327(B[327]),        // input wire [7 : 0] B_327
  .B_328(B[328]),        // input wire [7 : 0] B_328
  .B_329(B[329]),        // input wire [7 : 0] B_329
  .B_330(B[330]),        // input wire [7 : 0] B_330
  .B_331(B[331]),        // input wire [7 : 0] B_331
  .B_332(B[332]),        // input wire [7 : 0] B_332
  .B_333(B[333]),        // input wire [7 : 0] B_333
  .B_334(B[334]),        // input wire [7 : 0] B_334
  .B_335(B[335]),        // input wire [7 : 0] B_335
  .B_336(B[336]),        // input wire [7 : 0] B_336
  .B_337(B[337]),        // input wire [7 : 0] B_337
  .B_338(B[338]),        // input wire [7 : 0] B_338
  .B_339(B[339]),        // input wire [7 : 0] B_339
  .B_340(B[340]),        // input wire [7 : 0] B_340
  .B_341(B[341]),        // input wire [7 : 0] B_341
  .B_342(B[342]),        // input wire [7 : 0] B_342
  .B_343(B[343]),        // input wire [7 : 0] B_343
  .B_344(B[344]),        // input wire [7 : 0] B_344
  .B_345(B[345]),        // input wire [7 : 0] B_345
  .B_346(B[346]),        // input wire [7 : 0] B_346
  .B_347(B[347]),        // input wire [7 : 0] B_347
  .B_348(B[348]),        // input wire [7 : 0] B_348
  .B_349(B[349]),        // input wire [7 : 0] B_349
  .B_350(B[350]),        // input wire [7 : 0] B_350
  .B_351(B[351]),        // input wire [7 : 0] B_351
  .B_352(B[352]),        // input wire [7 : 0] B_352
  .B_353(B[353]),        // input wire [7 : 0] B_353
  .B_354(B[354]),        // input wire [7 : 0] B_354
  .B_355(B[355]),        // input wire [7 : 0] B_355
  .B_356(B[356]),        // input wire [7 : 0] B_356
  .B_357(B[357]),        // input wire [7 : 0] B_357
  .B_358(B[358]),        // input wire [7 : 0] B_358
  .B_359(B[359]),        // input wire [7 : 0] B_359
  .B_360(B[360]),        // input wire [7 : 0] B_360
  .B_361(B[361]),        // input wire [7 : 0] B_361
  .B_362(B[362]),        // input wire [7 : 0] B_362
  .B_363(B[363]),        // input wire [7 : 0] B_363
  .B_364(B[364]),        // input wire [7 : 0] B_364
  .B_365(B[365]),        // input wire [7 : 0] B_365
  .B_366(B[366]),        // input wire [7 : 0] B_366
  .B_367(B[367]),        // input wire [7 : 0] B_367
  .B_368(B[368]),        // input wire [7 : 0] B_368
  .B_369(B[369]),        // input wire [7 : 0] B_369
  .B_370(B[370]),        // input wire [7 : 0] B_370
  .B_371(B[371]),        // input wire [7 : 0] B_371
  .B_372(B[372]),        // input wire [7 : 0] B_372
  .B_373(B[373]),        // input wire [7 : 0] B_373
  .B_374(B[374]),        // input wire [7 : 0] B_374
  .B_375(B[375]),        // input wire [7 : 0] B_375
  .B_376(B[376]),        // input wire [7 : 0] B_376
  .B_377(B[377]),        // input wire [7 : 0] B_377
  .B_378(B[378]),        // input wire [7 : 0] B_378
  .B_379(B[379]),        // input wire [7 : 0] B_379
  .B_380(B[380]),        // input wire [7 : 0] B_380
  .B_381(B[381]),        // input wire [7 : 0] B_381
  .B_382(B[382]),        // input wire [7 : 0] B_382
  .B_383(B[383]),        // input wire [7 : 0] B_383
  .B_384(B[384]),        // input wire [7 : 0] B_384
  .B_385(B[385]),        // input wire [7 : 0] B_385
  .B_386(B[386]),        // input wire [7 : 0] B_386
  .B_387(B[387]),        // input wire [7 : 0] B_387
  .B_388(B[388]),        // input wire [7 : 0] B_388
  .B_389(B[389]),        // input wire [7 : 0] B_389
  .B_390(B[390]),        // input wire [7 : 0] B_390
  .B_391(B[391]),        // input wire [7 : 0] B_391
  .B_392(B[392]),        // input wire [7 : 0] B_392
  .B_393(B[393]),        // input wire [7 : 0] B_393
  .B_394(B[394]),        // input wire [7 : 0] B_394
  .B_395(B[395]),        // input wire [7 : 0] B_395
  .B_396(B[396]),        // input wire [7 : 0] B_396
  .B_397(B[397]),        // input wire [7 : 0] B_397
  .B_398(B[398]),        // input wire [7 : 0] B_398
  .B_399(B[399]),        // input wire [7 : 0] B_399
  .B_400(B[400]),        // input wire [7 : 0] B_400
  .B_401(B[401]),        // input wire [7 : 0] B_401
  .B_402(B[402]),        // input wire [7 : 0] B_402
  .B_403(B[403]),        // input wire [7 : 0] B_403
  .B_404(B[404]),        // input wire [7 : 0] B_404
  .B_405(B[405]),        // input wire [7 : 0] B_405
  .B_406(B[406]),        // input wire [7 : 0] B_406
  .B_407(B[407]),        // input wire [7 : 0] B_407
  .B_408(B[408]),        // input wire [7 : 0] B_408
  .B_409(B[409]),        // input wire [7 : 0] B_409
  .B_410(B[410]),        // input wire [7 : 0] B_410
  .B_411(B[411]),        // input wire [7 : 0] B_411
  .B_412(B[412]),        // input wire [7 : 0] B_412
  .B_413(B[413]),        // input wire [7 : 0] B_413
  .B_414(B[414]),        // input wire [7 : 0] B_414
  .B_415(B[415]),        // input wire [7 : 0] B_415
  .B_416(B[416]),        // input wire [7 : 0] B_416
  .B_417(B[417]),        // input wire [7 : 0] B_417
  .B_418(B[418]),        // input wire [7 : 0] B_418
  .B_419(B[419]),        // input wire [7 : 0] B_419
  .B_420(B[420]),        // input wire [7 : 0] B_420
  .B_421(B[421]),        // input wire [7 : 0] B_421
  .B_422(B[422]),        // input wire [7 : 0] B_422
  .B_423(B[423]),        // input wire [7 : 0] B_423
  .B_424(B[424]),        // input wire [7 : 0] B_424
  .B_425(B[425]),        // input wire [7 : 0] B_425
  .B_426(B[426]),        // input wire [7 : 0] B_426
  .B_427(B[427]),        // input wire [7 : 0] B_427
  .B_428(B[428]),        // input wire [7 : 0] B_428
  .B_429(B[429]),        // input wire [7 : 0] B_429
  .B_430(B[430]),        // input wire [7 : 0] B_430
  .B_431(B[431]),        // input wire [7 : 0] B_431
  .B_432(B[432]),        // input wire [7 : 0] B_432
  .B_433(B[433]),        // input wire [7 : 0] B_433
  .B_434(B[434]),        // input wire [7 : 0] B_434
  .B_435(B[435]),        // input wire [7 : 0] B_435
  .B_436(B[436]),        // input wire [7 : 0] B_436
  .B_437(B[437]),        // input wire [7 : 0] B_437
  .B_438(B[438]),        // input wire [7 : 0] B_438
  .B_439(B[439]),        // input wire [7 : 0] B_439
  .B_440(B[440]),        // input wire [7 : 0] B_440
  .B_441(B[441]),        // input wire [7 : 0] B_441
  .B_442(B[442]),        // input wire [7 : 0] B_442
  .B_443(B[443]),        // input wire [7 : 0] B_443
  .B_444(B[444]),        // input wire [7 : 0] B_444
  .B_445(B[445]),        // input wire [7 : 0] B_445
  .B_446(B[446]),        // input wire [7 : 0] B_446
  .B_447(B[447]),        // input wire [7 : 0] B_447
  .B_448(B[448]),        // input wire [7 : 0] B_448
  .B_449(B[449]),        // input wire [7 : 0] B_449
  .B_450(B[450]),        // input wire [7 : 0] B_450
  .B_451(B[451]),        // input wire [7 : 0] B_451
  .B_452(B[452]),        // input wire [7 : 0] B_452
  .B_453(B[453]),        // input wire [7 : 0] B_453
  .B_454(B[454]),        // input wire [7 : 0] B_454
  .B_455(B[455]),        // input wire [7 : 0] B_455
  .B_456(B[456]),        // input wire [7 : 0] B_456
  .B_457(B[457]),        // input wire [7 : 0] B_457
  .B_458(B[458]),        // input wire [7 : 0] B_458
  .B_459(B[459]),        // input wire [7 : 0] B_459
  .B_460(B[460]),        // input wire [7 : 0] B_460
  .B_461(B[461]),        // input wire [7 : 0] B_461
  .B_462(B[462]),        // input wire [7 : 0] B_462
  .B_463(B[463]),        // input wire [7 : 0] B_463
  .B_464(B[464]),        // input wire [7 : 0] B_464
  .B_465(B[465]),        // input wire [7 : 0] B_465
  .B_466(B[466]),        // input wire [7 : 0] B_466
  .B_467(B[467]),        // input wire [7 : 0] B_467
  .B_468(B[468]),        // input wire [7 : 0] B_468
  .B_469(B[469]),        // input wire [7 : 0] B_469
  .B_470(B[470]),        // input wire [7 : 0] B_470
  .B_471(B[471]),        // input wire [7 : 0] B_471
  .B_472(B[472]),        // input wire [7 : 0] B_472
  .B_473(B[473]),        // input wire [7 : 0] B_473
  .B_474(B[474]),        // input wire [7 : 0] B_474
  .B_475(B[475]),        // input wire [7 : 0] B_475
  .B_476(B[476]),        // input wire [7 : 0] B_476
  .B_477(B[477]),        // input wire [7 : 0] B_477
  .B_478(B[478]),        // input wire [7 : 0] B_478
  .B_479(B[479]),        // input wire [7 : 0] B_479
  .B_480(B[480]),        // input wire [7 : 0] B_480
  .B_481(B[481]),        // input wire [7 : 0] B_481
  .B_482(B[482]),        // input wire [7 : 0] B_482
  .B_483(B[483]),        // input wire [7 : 0] B_483
  .B_484(B[484]),        // input wire [7 : 0] B_484
  .B_485(B[485]),        // input wire [7 : 0] B_485
  .B_486(B[486]),        // input wire [7 : 0] B_486
  .B_487(B[487]),        // input wire [7 : 0] B_487
  .B_488(B[488]),        // input wire [7 : 0] B_488
  .B_489(B[489]),        // input wire [7 : 0] B_489
  .B_490(B[490]),        // input wire [7 : 0] B_490
  .B_491(B[491]),        // input wire [7 : 0] B_491
  .B_492(B[492]),        // input wire [7 : 0] B_492
  .B_493(B[493]),        // input wire [7 : 0] B_493
  .B_494(B[494]),        // input wire [7 : 0] B_494
  .B_495(B[495]),        // input wire [7 : 0] B_495
  .B_496(B[496]),        // input wire [7 : 0] B_496
  .B_497(B[497]),        // input wire [7 : 0] B_497
  .B_498(B[498]),        // input wire [7 : 0] B_498
  .B_499(B[499]),        // input wire [7 : 0] B_499
  .B_500(B[500]),        // input wire [7 : 0] B_500
  .B_501(B[501]),        // input wire [7 : 0] B_501
  .B_502(B[502]),        // input wire [7 : 0] B_502
  .B_503(B[503]),        // input wire [7 : 0] B_503
  .B_504(B[504]),        // input wire [7 : 0] B_504
  .B_505(B[505]),        // input wire [7 : 0] B_505
  .B_506(B[506]),        // input wire [7 : 0] B_506
  .B_507(B[507]),        // input wire [7 : 0] B_507
  .B_508(B[508]),        // input wire [7 : 0] B_508
  .B_509(B[509]),        // input wire [7 : 0] B_509
  .B_510(B[510]),        // input wire [7 : 0] B_510
  .B_511(B[511]),        // input wire [7 : 0] B_511
  .B_512(B[512]),        // input wire [7 : 0] B_512
  .B_513(B[513]),        // input wire [7 : 0] B_513
  .B_514(B[514]),        // input wire [7 : 0] B_514
  .B_515(B[515]),        // input wire [7 : 0] B_515
  .B_516(B[516]),        // input wire [7 : 0] B_516
  .B_517(B[517]),        // input wire [7 : 0] B_517
  .B_518(B[518]),        // input wire [7 : 0] B_518
  .B_519(B[519]),        // input wire [7 : 0] B_519
  .B_520(B[520]),        // input wire [7 : 0] B_520
  .B_521(B[521]),        // input wire [7 : 0] B_521
  .B_522(B[522]),        // input wire [7 : 0] B_522
  .B_523(B[523]),        // input wire [7 : 0] B_523
  .B_524(B[524]),        // input wire [7 : 0] B_524
  .B_525(B[525]),        // input wire [7 : 0] B_525
  .B_526(B[526]),        // input wire [7 : 0] B_526
  .B_527(B[527]),        // input wire [7 : 0] B_527
  .B_528(B[528]),        // input wire [7 : 0] B_528
  .B_529(B[529]),        // input wire [7 : 0] B_529
  .B_530(B[530]),        // input wire [7 : 0] B_530
  .B_531(B[531]),        // input wire [7 : 0] B_531
  .B_532(B[532]),        // input wire [7 : 0] B_532
  .B_533(B[533]),        // input wire [7 : 0] B_533
  .B_534(B[534]),        // input wire [7 : 0] B_534
  .B_535(B[535]),        // input wire [7 : 0] B_535
  .B_536(B[536]),        // input wire [7 : 0] B_536
  .B_537(B[537]),        // input wire [7 : 0] B_537
  .B_538(B[538]),        // input wire [7 : 0] B_538
  .B_539(B[539]),        // input wire [7 : 0] B_539
  .B_540(B[540]),        // input wire [7 : 0] B_540
  .B_541(B[541]),        // input wire [7 : 0] B_541
  .B_542(B[542]),        // input wire [7 : 0] B_542
  .B_543(B[543]),        // input wire [7 : 0] B_543
  .B_544(B[544]),        // input wire [7 : 0] B_544
  .B_545(B[545]),        // input wire [7 : 0] B_545
  .B_546(B[546]),        // input wire [7 : 0] B_546
  .B_547(B[547]),        // input wire [7 : 0] B_547
  .B_548(B[548]),        // input wire [7 : 0] B_548
  .B_549(B[549]),        // input wire [7 : 0] B_549
  .B_550(B[550]),        // input wire [7 : 0] B_550
  .B_551(B[551]),        // input wire [7 : 0] B_551
  .B_552(B[552]),        // input wire [7 : 0] B_552
  .B_553(B[553]),        // input wire [7 : 0] B_553
  .B_554(B[554]),        // input wire [7 : 0] B_554
  .B_555(B[555]),        // input wire [7 : 0] B_555
  .B_556(B[556]),        // input wire [7 : 0] B_556
  .B_557(B[557]),        // input wire [7 : 0] B_557
  .B_558(B[558]),        // input wire [7 : 0] B_558
  .B_559(B[559]),        // input wire [7 : 0] B_559
  .B_560(B[560]),        // input wire [7 : 0] B_560
  .B_561(B[561]),        // input wire [7 : 0] B_561
  .B_562(B[562]),        // input wire [7 : 0] B_562
  .B_563(B[563]),        // input wire [7 : 0] B_563
  .B_564(B[564]),        // input wire [7 : 0] B_564
  .B_565(B[565]),        // input wire [7 : 0] B_565
  .B_566(B[566]),        // input wire [7 : 0] B_566
  .B_567(B[567]),        // input wire [7 : 0] B_567
  .B_568(B[568]),        // input wire [7 : 0] B_568
  .B_569(B[569]),        // input wire [7 : 0] B_569
  .B_570(B[570]),        // input wire [7 : 0] B_570
  .B_571(B[571]),        // input wire [7 : 0] B_571
  .B_572(B[572]),        // input wire [7 : 0] B_572
  .B_573(B[573]),        // input wire [7 : 0] B_573
  .B_574(B[574]),        // input wire [7 : 0] B_574
  .B_575(B[575]),        // input wire [7 : 0] B_575
  .B_576(B[576]),        // input wire [7 : 0] B_576
  .B_577(B[577]),        // input wire [7 : 0] B_577
  .B_578(B[578]),        // input wire [7 : 0] B_578
  .B_579(B[579]),        // input wire [7 : 0] B_579
  .B_580(B[580]),        // input wire [7 : 0] B_580
  .B_581(B[581]),        // input wire [7 : 0] B_581
  .B_582(B[582]),        // input wire [7 : 0] B_582
  .B_583(B[583]),        // input wire [7 : 0] B_583
  .B_584(B[584]),        // input wire [7 : 0] B_584
  .B_585(B[585]),        // input wire [7 : 0] B_585
  .B_586(B[586]),        // input wire [7 : 0] B_586
  .B_587(B[587]),        // input wire [7 : 0] B_587
  .B_588(B[588]),        // input wire [7 : 0] B_588
  .B_589(B[589]),        // input wire [7 : 0] B_589
  .B_590(B[590]),        // input wire [7 : 0] B_590
  .B_591(B[591]),        // input wire [7 : 0] B_591
  .B_592(B[592]),        // input wire [7 : 0] B_592
  .B_593(B[593]),        // input wire [7 : 0] B_593
  .B_594(B[594]),        // input wire [7 : 0] B_594
  .B_595(B[595]),        // input wire [7 : 0] B_595
  .B_596(B[596]),        // input wire [7 : 0] B_596
  .B_597(B[597]),        // input wire [7 : 0] B_597
  .B_598(B[598]),        // input wire [7 : 0] B_598
  .B_599(B[599]),        // input wire [7 : 0] B_599
  .B_600(B[600]),        // input wire [7 : 0] B_600
  .B_601(B[601]),        // input wire [7 : 0] B_601
  .B_602(B[602]),        // input wire [7 : 0] B_602
  .B_603(B[603]),        // input wire [7 : 0] B_603
  .B_604(B[604]),        // input wire [7 : 0] B_604
  .B_605(B[605]),        // input wire [7 : 0] B_605
  .B_606(B[606]),        // input wire [7 : 0] B_606
  .B_607(B[607]),        // input wire [7 : 0] B_607
  .B_608(B[608]),        // input wire [7 : 0] B_608
  .B_609(B[609]),        // input wire [7 : 0] B_609
  .B_610(B[610]),        // input wire [7 : 0] B_610
  .B_611(B[611]),        // input wire [7 : 0] B_611
  .B_612(B[612]),        // input wire [7 : 0] B_612
  .B_613(B[613]),        // input wire [7 : 0] B_613
  .B_614(B[614]),        // input wire [7 : 0] B_614
  .B_615(B[615]),        // input wire [7 : 0] B_615
  .B_616(B[616]),        // input wire [7 : 0] B_616
  .B_617(B[617]),        // input wire [7 : 0] B_617
  .B_618(B[618]),        // input wire [7 : 0] B_618
  .B_619(B[619]),        // input wire [7 : 0] B_619
  .B_620(B[620]),        // input wire [7 : 0] B_620
  .B_621(B[621]),        // input wire [7 : 0] B_621
  .B_622(B[622]),        // input wire [7 : 0] B_622
  .B_623(B[623]),        // input wire [7 : 0] B_623
  .B_624(B[624]),        // input wire [7 : 0] B_624
  .B_625(B[625]),        // input wire [7 : 0] B_625
  .B_626(B[626]),        // input wire [7 : 0] B_626
  .B_627(B[627]),        // input wire [7 : 0] B_627
  .B_628(B[628]),        // input wire [7 : 0] B_628
  .B_629(B[629]),        // input wire [7 : 0] B_629
  .B_630(B[630]),        // input wire [7 : 0] B_630
  .B_631(B[631]),        // input wire [7 : 0] B_631
  .B_632(B[632]),        // input wire [7 : 0] B_632
  .B_633(B[633]),        // input wire [7 : 0] B_633
  .B_634(B[634]),        // input wire [7 : 0] B_634
  .B_635(B[635]),        // input wire [7 : 0] B_635
  .B_636(B[636]),        // input wire [7 : 0] B_636
  .B_637(B[637]),        // input wire [7 : 0] B_637
  .B_638(B[638]),        // input wire [7 : 0] B_638
  .B_639(B[639]),        // input wire [7 : 0] B_639
  .B_640(B[640]),        // input wire [7 : 0] B_640
  .B_641(B[641]),        // input wire [7 : 0] B_641
  .B_642(B[642]),        // input wire [7 : 0] B_642
  .B_643(B[643]),        // input wire [7 : 0] B_643
  .B_644(B[644]),        // input wire [7 : 0] B_644
  .B_645(B[645]),        // input wire [7 : 0] B_645
  .B_646(B[646]),        // input wire [7 : 0] B_646
  .B_647(B[647]),        // input wire [7 : 0] B_647
  .B_648(B[648]),        // input wire [7 : 0] B_648
  .B_649(B[649]),        // input wire [7 : 0] B_649
  .B_650(B[650]),        // input wire [7 : 0] B_650
  .B_651(B[651]),        // input wire [7 : 0] B_651
  .B_652(B[652]),        // input wire [7 : 0] B_652
  .B_653(B[653]),        // input wire [7 : 0] B_653
  .B_654(B[654]),        // input wire [7 : 0] B_654
  .B_655(B[655]),        // input wire [7 : 0] B_655
  .B_656(B[656]),        // input wire [7 : 0] B_656
  .B_657(B[657]),        // input wire [7 : 0] B_657
  .B_658(B[658]),        // input wire [7 : 0] B_658
  .B_659(B[659]),        // input wire [7 : 0] B_659
  .B_660(B[660]),        // input wire [7 : 0] B_660
  .B_661(B[661]),        // input wire [7 : 0] B_661
  .B_662(B[662]),        // input wire [7 : 0] B_662
  .B_663(B[663]),        // input wire [7 : 0] B_663
  .B_664(B[664]),        // input wire [7 : 0] B_664
  .B_665(B[665]),        // input wire [7 : 0] B_665
  .B_666(B[666]),        // input wire [7 : 0] B_666
  .B_667(B[667]),        // input wire [7 : 0] B_667
  .B_668(B[668]),        // input wire [7 : 0] B_668
  .B_669(B[669]),        // input wire [7 : 0] B_669
  .B_670(B[670]),        // input wire [7 : 0] B_670
  .B_671(B[671]),        // input wire [7 : 0] B_671
  .B_672(B[672]),        // input wire [7 : 0] B_672
  .B_673(B[673]),        // input wire [7 : 0] B_673
  .B_674(B[674]),        // input wire [7 : 0] B_674
  .B_675(B[675]),        // input wire [7 : 0] B_675
  .B_676(B[676]),        // input wire [7 : 0] B_676
  .B_677(B[677]),        // input wire [7 : 0] B_677
  .B_678(B[678]),        // input wire [7 : 0] B_678
  .B_679(B[679]),        // input wire [7 : 0] B_679
  .B_680(B[680]),        // input wire [7 : 0] B_680
  .B_681(B[681]),        // input wire [7 : 0] B_681
  .B_682(B[682]),        // input wire [7 : 0] B_682
  .B_683(B[683]),        // input wire [7 : 0] B_683
  .B_684(B[684]),        // input wire [7 : 0] B_684
  .B_685(B[685]),        // input wire [7 : 0] B_685
  .B_686(B[686]),        // input wire [7 : 0] B_686
  .B_687(B[687]),        // input wire [7 : 0] B_687
  .B_688(B[688]),        // input wire [7 : 0] B_688
  .B_689(B[689]),        // input wire [7 : 0] B_689
  .B_690(B[690]),        // input wire [7 : 0] B_690
  .B_691(B[691]),        // input wire [7 : 0] B_691
  .B_692(B[692]),        // input wire [7 : 0] B_692
  .B_693(B[693]),        // input wire [7 : 0] B_693
  .B_694(B[694]),        // input wire [7 : 0] B_694
  .B_695(B[695]),        // input wire [7 : 0] B_695
  .B_696(B[696]),        // input wire [7 : 0] B_696
  .B_697(B[697]),        // input wire [7 : 0] B_697
  .B_698(B[698]),        // input wire [7 : 0] B_698
  .B_699(B[699]),        // input wire [7 : 0] B_699
  .B_700(B[700]),        // input wire [7 : 0] B_700
  .B_701(B[701]),        // input wire [7 : 0] B_701
  .B_702(B[702]),        // input wire [7 : 0] B_702
  .B_703(B[703]),        // input wire [7 : 0] B_703
  .B_704(B[704]),        // input wire [7 : 0] B_704
  .B_705(B[705]),        // input wire [7 : 0] B_705
  .B_706(B[706]),        // input wire [7 : 0] B_706
  .B_707(B[707]),        // input wire [7 : 0] B_707
  .B_708(B[708]),        // input wire [7 : 0] B_708
  .B_709(B[709]),        // input wire [7 : 0] B_709
  .B_710(B[710]),        // input wire [7 : 0] B_710
  .B_711(B[711]),        // input wire [7 : 0] B_711
  .B_712(B[712]),        // input wire [7 : 0] B_712
  .B_713(B[713]),        // input wire [7 : 0] B_713
  .B_714(B[714]),        // input wire [7 : 0] B_714
  .B_715(B[715]),        // input wire [7 : 0] B_715
  .B_716(B[716]),        // input wire [7 : 0] B_716
  .B_717(B[717]),        // input wire [7 : 0] B_717
  .B_718(B[718]),        // input wire [7 : 0] B_718
  .B_719(B[719]),        // input wire [7 : 0] B_719
  .B_720(B[720]),        // input wire [7 : 0] B_720
  .B_721(B[721]),        // input wire [7 : 0] B_721
  .B_722(B[722]),        // input wire [7 : 0] B_722
  .B_723(B[723]),        // input wire [7 : 0] B_723
  .B_724(B[724]),        // input wire [7 : 0] B_724
  .B_725(B[725]),        // input wire [7 : 0] B_725
  .B_726(B[726]),        // input wire [7 : 0] B_726
  .B_727(B[727]),        // input wire [7 : 0] B_727
  .B_728(B[728]),        // input wire [7 : 0] B_728
  .B_729(B[729]),        // input wire [7 : 0] B_729
  .B_730(B[730]),        // input wire [7 : 0] B_730
  .B_731(B[731]),        // input wire [7 : 0] B_731
  .B_732(B[732]),        // input wire [7 : 0] B_732
  .B_733(B[733]),        // input wire [7 : 0] B_733
  .B_734(B[734]),        // input wire [7 : 0] B_734
  .B_735(B[735]),        // input wire [7 : 0] B_735
  .B_736(B[736]),        // input wire [7 : 0] B_736
  .B_737(B[737]),        // input wire [7 : 0] B_737
  .B_738(B[738]),        // input wire [7 : 0] B_738
  .B_739(B[739]),        // input wire [7 : 0] B_739
  .B_740(B[740]),        // input wire [7 : 0] B_740
  .B_741(B[741]),        // input wire [7 : 0] B_741
  .B_742(B[742]),        // input wire [7 : 0] B_742
  .B_743(B[743]),        // input wire [7 : 0] B_743
  .B_744(B[744]),        // input wire [7 : 0] B_744
  .B_745(B[745]),        // input wire [7 : 0] B_745
  .B_746(B[746]),        // input wire [7 : 0] B_746
  .B_747(B[747]),        // input wire [7 : 0] B_747
  .B_748(B[748]),        // input wire [7 : 0] B_748
  .B_749(B[749]),        // input wire [7 : 0] B_749
  .B_750(B[750]),        // input wire [7 : 0] B_750
  .B_751(B[751]),        // input wire [7 : 0] B_751
  .B_752(B[752]),        // input wire [7 : 0] B_752
  .B_753(B[753]),        // input wire [7 : 0] B_753
  .B_754(B[754]),        // input wire [7 : 0] B_754
  .B_755(B[755]),        // input wire [7 : 0] B_755
  .B_756(B[756]),        // input wire [7 : 0] B_756
  .B_757(B[757]),        // input wire [7 : 0] B_757
  .B_758(B[758]),        // input wire [7 : 0] B_758
  .B_759(B[759]),        // input wire [7 : 0] B_759
  .B_760(B[760]),        // input wire [7 : 0] B_760
  .B_761(B[761]),        // input wire [7 : 0] B_761
  .B_762(B[762]),        // input wire [7 : 0] B_762
  .B_763(B[763]),        // input wire [7 : 0] B_763
  .B_764(B[764]),        // input wire [7 : 0] B_764
  .B_765(B[765]),        // input wire [7 : 0] B_765
  .B_766(B[766]),        // input wire [7 : 0] B_766
  .B_767(B[767]),        // input wire [7 : 0] B_767
  .B_768(B[768]),        // input wire [7 : 0] B_768
  .B_769(B[769]),        // input wire [7 : 0] B_769
  .B_770(B[770]),        // input wire [7 : 0] B_770
  .B_771(B[771]),        // input wire [7 : 0] B_771
  .B_772(B[772]),        // input wire [7 : 0] B_772
  .B_773(B[773]),        // input wire [7 : 0] B_773
  .B_774(B[774]),        // input wire [7 : 0] B_774
  .B_775(B[775]),        // input wire [7 : 0] B_775
  .B_776(B[776]),        // input wire [7 : 0] B_776
  .B_777(B[777]),        // input wire [7 : 0] B_777
  .B_778(B[778]),        // input wire [7 : 0] B_778
  .B_779(B[779]),        // input wire [7 : 0] B_779
  .B_780(B[780]),        // input wire [7 : 0] B_780
  .B_781(B[781]),        // input wire [7 : 0] B_781
  .B_782(B[782]),        // input wire [7 : 0] B_782
  .B_783(B[783]),        // input wire [7 : 0] B_783
  .B_784(B[784]),        // input wire [7 : 0] B_784
  .B_785(B[785]),        // input wire [7 : 0] B_785
  .B_786(B[786]),        // input wire [7 : 0] B_786
  .B_787(B[787]),        // input wire [7 : 0] B_787
  .B_788(B[788]),        // input wire [7 : 0] B_788
  .B_789(B[789]),        // input wire [7 : 0] B_789
  .B_790(B[790]),        // input wire [7 : 0] B_790
  .B_791(B[791]),        // input wire [7 : 0] B_791
  .B_792(B[792]),        // input wire [7 : 0] B_792
  .B_793(B[793]),        // input wire [7 : 0] B_793
  .B_794(B[794]),        // input wire [7 : 0] B_794
  .B_795(B[795]),        // input wire [7 : 0] B_795
  .B_796(B[796]),        // input wire [7 : 0] B_796
  .B_797(B[797]),        // input wire [7 : 0] B_797
  .B_798(B[798]),        // input wire [7 : 0] B_798
  .B_799(B[799]),        // input wire [7 : 0] B_799
  .B_800(B[800]),        // input wire [7 : 0] B_800
  .B_801(B[801]),        // input wire [7 : 0] B_801
  .B_802(B[802]),        // input wire [7 : 0] B_802
  .B_803(B[803]),        // input wire [7 : 0] B_803
  .B_804(B[804]),        // input wire [7 : 0] B_804
  .B_805(B[805]),        // input wire [7 : 0] B_805
  .B_806(B[806]),        // input wire [7 : 0] B_806
  .B_807(B[807]),        // input wire [7 : 0] B_807
  .B_808(B[808]),        // input wire [7 : 0] B_808
  .B_809(B[809]),        // input wire [7 : 0] B_809
  .B_810(B[810]),        // input wire [7 : 0] B_810
  .B_811(B[811]),        // input wire [7 : 0] B_811
  .B_812(B[812]),        // input wire [7 : 0] B_812
  .B_813(B[813]),        // input wire [7 : 0] B_813
  .B_814(B[814]),        // input wire [7 : 0] B_814
  .B_815(B[815]),        // input wire [7 : 0] B_815
  .B_816(B[816]),        // input wire [7 : 0] B_816
  .B_817(B[817]),        // input wire [7 : 0] B_817
  .B_818(B[818]),        // input wire [7 : 0] B_818
  .B_819(B[819]),        // input wire [7 : 0] B_819
  .B_820(B[820]),        // input wire [7 : 0] B_820
  .B_821(B[821]),        // input wire [7 : 0] B_821
  .B_822(B[822]),        // input wire [7 : 0] B_822
  .B_823(B[823]),        // input wire [7 : 0] B_823
  .B_824(B[824]),        // input wire [7 : 0] B_824
  .B_825(B[825]),        // input wire [7 : 0] B_825
  .B_826(B[826]),        // input wire [7 : 0] B_826
  .B_827(B[827]),        // input wire [7 : 0] B_827
  .B_828(B[828]),        // input wire [7 : 0] B_828
  .B_829(B[829]),        // input wire [7 : 0] B_829
  .B_830(B[830]),        // input wire [7 : 0] B_830
  .B_831(B[831]),        // input wire [7 : 0] B_831
  .B_832(B[832]),        // input wire [7 : 0] B_832
  .B_833(B[833]),        // input wire [7 : 0] B_833
  .B_834(B[834]),        // input wire [7 : 0] B_834
  .B_835(B[835]),        // input wire [7 : 0] B_835
  .B_836(B[836]),        // input wire [7 : 0] B_836
  .B_837(B[837]),        // input wire [7 : 0] B_837
  .B_838(B[838]),        // input wire [7 : 0] B_838
  .B_839(B[839]),        // input wire [7 : 0] B_839
  .B_840(B[840]),        // input wire [7 : 0] B_840
  .B_841(B[841]),        // input wire [7 : 0] B_841
  .B_842(B[842]),        // input wire [7 : 0] B_842
  .B_843(B[843]),        // input wire [7 : 0] B_843
  .B_844(B[844]),        // input wire [7 : 0] B_844
  .B_845(B[845]),        // input wire [7 : 0] B_845
  .B_846(B[846]),        // input wire [7 : 0] B_846
  .B_847(B[847]),        // input wire [7 : 0] B_847
  .B_848(B[848]),        // input wire [7 : 0] B_848
  .B_849(B[849]),        // input wire [7 : 0] B_849
  .B_850(B[850]),        // input wire [7 : 0] B_850
  .B_851(B[851]),        // input wire [7 : 0] B_851
  .B_852(B[852]),        // input wire [7 : 0] B_852
  .B_853(B[853]),        // input wire [7 : 0] B_853
  .B_854(B[854]),        // input wire [7 : 0] B_854
  .B_855(B[855]),        // input wire [7 : 0] B_855
  .B_856(B[856]),        // input wire [7 : 0] B_856
  .B_857(B[857]),        // input wire [7 : 0] B_857
  .B_858(B[858]),        // input wire [7 : 0] B_858
  .B_859(B[859]),        // input wire [7 : 0] B_859
  .B_860(B[860]),        // input wire [7 : 0] B_860
  .B_861(B[861]),        // input wire [7 : 0] B_861
  .B_862(B[862]),        // input wire [7 : 0] B_862
  .B_863(B[863]),        // input wire [7 : 0] B_863
  .B_864(B[864]),        // input wire [7 : 0] B_864
  .B_865(B[865]),        // input wire [7 : 0] B_865
  .B_866(B[866]),        // input wire [7 : 0] B_866
  .B_867(B[867]),        // input wire [7 : 0] B_867
  .B_868(B[868]),        // input wire [7 : 0] B_868
  .B_869(B[869]),        // input wire [7 : 0] B_869
  .B_870(B[870]),        // input wire [7 : 0] B_870
  .B_871(B[871]),        // input wire [7 : 0] B_871
  .B_872(B[872]),        // input wire [7 : 0] B_872
  .B_873(B[873]),        // input wire [7 : 0] B_873
  .B_874(B[874]),        // input wire [7 : 0] B_874
  .B_875(B[875]),        // input wire [7 : 0] B_875
  .B_876(B[876]),        // input wire [7 : 0] B_876
  .B_877(B[877]),        // input wire [7 : 0] B_877
  .B_878(B[878]),        // input wire [7 : 0] B_878
  .B_879(B[879]),        // input wire [7 : 0] B_879
  .B_880(B[880]),        // input wire [7 : 0] B_880
  .B_881(B[881]),        // input wire [7 : 0] B_881
  .B_882(B[882]),        // input wire [7 : 0] B_882
  .B_883(B[883]),        // input wire [7 : 0] B_883
  .B_884(B[884]),        // input wire [7 : 0] B_884
  .B_885(B[885]),        // input wire [7 : 0] B_885
  .B_886(B[886]),        // input wire [7 : 0] B_886
  .B_887(B[887]),        // input wire [7 : 0] B_887
  .B_888(B[888]),        // input wire [7 : 0] B_888
  .B_889(B[889]),        // input wire [7 : 0] B_889
  .B_890(B[890]),        // input wire [7 : 0] B_890
  .B_891(B[891]),        // input wire [7 : 0] B_891
  .B_892(B[892]),        // input wire [7 : 0] B_892
  .B_893(B[893]),        // input wire [7 : 0] B_893
  .B_894(B[894]),        // input wire [7 : 0] B_894
  .B_895(B[895]),        // input wire [7 : 0] B_895
  .B_896(B[896]),        // input wire [7 : 0] B_896
  .B_897(B[897]),        // input wire [7 : 0] B_897
  .B_898(B[898]),        // input wire [7 : 0] B_898
  .B_899(B[899]),        // input wire [7 : 0] B_899
  .B_900(B[900]),        // input wire [7 : 0] B_900
  .B_901(B[901]),        // input wire [7 : 0] B_901
  .B_902(B[902]),        // input wire [7 : 0] B_902
  .B_903(B[903]),        // input wire [7 : 0] B_903
  .B_904(B[904]),        // input wire [7 : 0] B_904
  .B_905(B[905]),        // input wire [7 : 0] B_905
  .B_906(B[906]),        // input wire [7 : 0] B_906
  .B_907(B[907]),        // input wire [7 : 0] B_907
  .B_908(B[908]),        // input wire [7 : 0] B_908
  .B_909(B[909]),        // input wire [7 : 0] B_909
  .B_910(B[910]),        // input wire [7 : 0] B_910
  .B_911(B[911]),        // input wire [7 : 0] B_911
  .B_912(B[912]),        // input wire [7 : 0] B_912
  .B_913(B[913]),        // input wire [7 : 0] B_913
  .B_914(B[914]),        // input wire [7 : 0] B_914
  .B_915(B[915]),        // input wire [7 : 0] B_915
  .B_916(B[916]),        // input wire [7 : 0] B_916
  .B_917(B[917]),        // input wire [7 : 0] B_917
  .B_918(B[918]),        // input wire [7 : 0] B_918
  .B_919(B[919]),        // input wire [7 : 0] B_919
  .B_920(B[920]),        // input wire [7 : 0] B_920
  .B_921(B[921]),        // input wire [7 : 0] B_921
  .B_922(B[922]),        // input wire [7 : 0] B_922
  .B_923(B[923]),        // input wire [7 : 0] B_923
  .B_924(B[924]),        // input wire [7 : 0] B_924
  .B_925(B[925]),        // input wire [7 : 0] B_925
  .B_926(B[926]),        // input wire [7 : 0] B_926
  .B_927(B[927]),        // input wire [7 : 0] B_927
  .B_928(B[928]),        // input wire [7 : 0] B_928
  .B_929(B[929]),        // input wire [7 : 0] B_929
  .B_930(B[930]),        // input wire [7 : 0] B_930
  .B_931(B[931]),        // input wire [7 : 0] B_931
  .B_932(B[932]),        // input wire [7 : 0] B_932
  .B_933(B[933]),        // input wire [7 : 0] B_933
  .B_934(B[934]),        // input wire [7 : 0] B_934
  .B_935(B[935]),        // input wire [7 : 0] B_935
  .B_936(B[936]),        // input wire [7 : 0] B_936
  .B_937(B[937]),        // input wire [7 : 0] B_937
  .B_938(B[938]),        // input wire [7 : 0] B_938
  .B_939(B[939]),        // input wire [7 : 0] B_939
  .B_940(B[940]),        // input wire [7 : 0] B_940
  .B_941(B[941]),        // input wire [7 : 0] B_941
  .B_942(B[942]),        // input wire [7 : 0] B_942
  .B_943(B[943]),        // input wire [7 : 0] B_943
  .B_944(B[944]),        // input wire [7 : 0] B_944
  .B_945(B[945]),        // input wire [7 : 0] B_945
  .B_946(B[946]),        // input wire [7 : 0] B_946
  .B_947(B[947]),        // input wire [7 : 0] B_947
  .B_948(B[948]),        // input wire [7 : 0] B_948
  .B_949(B[949]),        // input wire [7 : 0] B_949
  .B_950(B[950]),        // input wire [7 : 0] B_950
  .B_951(B[951]),        // input wire [7 : 0] B_951
  .B_952(B[952]),        // input wire [7 : 0] B_952
  .B_953(B[953]),        // input wire [7 : 0] B_953
  .B_954(B[954]),        // input wire [7 : 0] B_954
  .B_955(B[955]),        // input wire [7 : 0] B_955
  .B_956(B[956]),        // input wire [7 : 0] B_956
  .B_957(B[957]),        // input wire [7 : 0] B_957
  .B_958(B[958]),        // input wire [7 : 0] B_958
  .B_959(B[959]),        // input wire [7 : 0] B_959
  .B_960(B[960]),        // input wire [7 : 0] B_960
  .B_961(B[961]),        // input wire [7 : 0] B_961
  .B_962(B[962]),        // input wire [7 : 0] B_962
  .B_963(B[963]),        // input wire [7 : 0] B_963
  .B_964(B[964]),        // input wire [7 : 0] B_964
  .B_965(B[965]),        // input wire [7 : 0] B_965
  .B_966(B[966]),        // input wire [7 : 0] B_966
  .B_967(B[967]),        // input wire [7 : 0] B_967
  .B_968(B[968]),        // input wire [7 : 0] B_968
  .B_969(B[969]),        // input wire [7 : 0] B_969
  .B_970(B[970]),        // input wire [7 : 0] B_970
  .B_971(B[971]),        // input wire [7 : 0] B_971
  .B_972(B[972]),        // input wire [7 : 0] B_972
  .B_973(B[973]),        // input wire [7 : 0] B_973
  .B_974(B[974]),        // input wire [7 : 0] B_974
  .B_975(B[975]),        // input wire [7 : 0] B_975
  .B_976(B[976]),        // input wire [7 : 0] B_976
  .B_977(B[977]),        // input wire [7 : 0] B_977
  .B_978(B[978]),        // input wire [7 : 0] B_978
  .B_979(B[979]),        // input wire [7 : 0] B_979
  .B_980(B[980]),        // input wire [7 : 0] B_980
  .B_981(B[981]),        // input wire [7 : 0] B_981
  .B_982(B[982]),        // input wire [7 : 0] B_982
  .B_983(B[983]),        // input wire [7 : 0] B_983
  .B_984(B[984]),        // input wire [7 : 0] B_984
  .B_985(B[985]),        // input wire [7 : 0] B_985
  .B_986(B[986]),        // input wire [7 : 0] B_986
  .B_987(B[987]),        // input wire [7 : 0] B_987
  .B_988(B[988]),        // input wire [7 : 0] B_988
  .B_989(B[989]),        // input wire [7 : 0] B_989
  .B_990(B[990]),        // input wire [7 : 0] B_990
  .B_991(B[991]),        // input wire [7 : 0] B_991
  .B_992(B[992]),        // input wire [7 : 0] B_992
  .B_993(B[993]),        // input wire [7 : 0] B_993
  .B_994(B[994]),        // input wire [7 : 0] B_994
  .B_995(B[995]),        // input wire [7 : 0] B_995
  .B_996(B[996]),        // input wire [7 : 0] B_996
  .B_997(B[997]),        // input wire [7 : 0] B_997
  .B_998(B[998]),        // input wire [7 : 0] B_998
  .B_999(B[999]),        // input wire [7 : 0] B_999
  .B_1000(B[1000]),      // input wire [7 : 0] B_1000
  .B_1001(B[1001]),      // input wire [7 : 0] B_1001
  .B_1002(B[1002]),      // input wire [7 : 0] B_1002
  .B_1003(B[1003]),      // input wire [7 : 0] B_1003
  .B_1004(B[1004]),      // input wire [7 : 0] B_1004
  .B_1005(B[1005]),      // input wire [7 : 0] B_1005
  .B_1006(B[1006]),      // input wire [7 : 0] B_1006
  .B_1007(B[1007]),      // input wire [7 : 0] B_1007
  .B_1008(B[1008]),      // input wire [7 : 0] B_1008
  .B_1009(B[1009]),      // input wire [7 : 0] B_1009
  .B_1010(B[1010]),      // input wire [7 : 0] B_1010
  .B_1011(B[1011]),      // input wire [7 : 0] B_1011
  .B_1012(B[1012]),      // input wire [7 : 0] B_1012
  .B_1013(B[1013]),      // input wire [7 : 0] B_1013
  .B_1014(B[1014]),      // input wire [7 : 0] B_1014
  .B_1015(B[1015]),      // input wire [7 : 0] B_1015
  .B_1016(B[1016]),      // input wire [7 : 0] B_1016
  .B_1017(B[1017]),      // input wire [7 : 0] B_1017
  .B_1018(B[1018]),      // input wire [7 : 0] B_1018
  .B_1019(B[1019]),      // input wire [7 : 0] B_1019
  .B_1020(B[1020]),      // input wire [7 : 0] B_1020
  .B_1021(B[1021]),      // input wire [7 : 0] B_1021
  .B_1022(B[1022]),      // input wire [7 : 0] B_1022
  .B_1023(B[1023]),      // input wire [7 : 0] B_1023
  .C(out)                // output wire [31 : 0] C
  );


endmodule
